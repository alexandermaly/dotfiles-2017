MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ��I�|��|��|�=���|�����|�is��|��|��|����|����n|�����|�����|�Rich�|�        PE  L �YU        � !    �     0�                               �                              �� G   �� x                            � ��  �#                            ض @              h                          .text   �                        `.rdata  �     �                @  @.data   ��   �  P   �             @  �.reloc  �"  �  0  @             @  B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �-w �����������U��W�}��xS�]V�u����u��y�^[_]� ���������� ��8��t�xu觴  ��t	�L  ��u3���  ��uø   ���������+ �� ������U��E�� t$��u��8�F4 ��u3�]��) �����]ø   ]�����������U���8V��H�QV�ҡ�8�H�U�AVR�Ѓ���^]� U���8V��H�QV�ҡ�8�U�H�E�IRj�PV�у���^]� ���������̡�8�P�BQ��Yø   @� ��������U��j�hd d�    PQV�  3�P�E�d�    ��u��8�H�QV�ҋ�8�Q�FP�B�E�    �Ћ�8�Q�F P�B�E��Ћ�8�Q�F0P�B�E��Ћ�8�Q�F@P�B�E��Ћ�8�Q�J�FPP�E��у��ƋM�d�    Y^��]����U��j�h� d�    PQV�  3�P�E�d�    ��u��8�H�A�VPR�E�   �Ћ�8�Q�J�F@P�E��ы�8�B�P�N0Q�E��ҡ�8�H�A�V R�E��Ћ�8�Q�J�FP�E� �ы�8�B�HV�E������у��M�d�    Y^��]����������������U��j�h!d�    P��dSV�  3�P�E�d�    �u�E�    ��8�P�Bdj�M�E�   ��h�#j�XhD�S�E��@ ��8�Q��jS�E�P�Bh�M�Ћ�8�Q�BV�Ѓ��}� �E�   �E�    ��  �M�U��
��/v��:r(��@v��[r��`v��{r��-t��_t
��.t��~ua��8�H�A�U�R�Ћ�8�Q�Rf�ÍM�PjQ�҃���8�P�B<���E��Ћ�8�Q�RLj�j��M�QP���ҍU���  �� ��8�Q�JuX�E�P�ы�8�B�Pj j��M�h�#Q�҃���8�P�B<���E��Ћ�8�Q�RLj�j��M�QP���ҍU��o  �E�P�ы�8�B�Pj j��M�h�#Q�҃���8�P�B<���E��Ћ�8�Q�RLj�j��M�QP���ҡ�8�H�A�U�R�E��Њ�����<	��v��7���0��8�Q�J�E�E�P��f�M��8�B�@�U�QjR�Ѓ���8�Q�B<���E��Ћ�8�Q�RLj�j��M�QP���ҡ�8�H�A�U�R�E����Ã�%  �yH���@<	��v��7���0��8�Q�J�E�P�ы�8�B�@f�ˍU�QjR�Ѓ���8�Q�B<���E��Ћ�8�Q�RLj�j��M�QP���ҍU���8�H�AR�E��ЋE�����;E�E��e����E��t	P�a< ����8�Q�J�EP�E� �у��ƋM�d�    Y^[��]���U��j�hM!d�    PQV�  3�P�E�d�    h�#j}hD�j�y< �����u����E�    t���o3 ��#���3�Ph'  �E�������8�$ ��Pj j h'  ��# ��Phi� �|5 ���M�d�    Y^��]����������U��j�h�!d�    PQV�  3�P�E�d�    �E�    ��8�H�u�QV�E�    �ҡ�8�H�U�AVR�Ѓ���8�Q�B<���E�    �E�   �Ћ�8�Q�M�RLj�j�QP���ҋƋM�d�    Y^��]����������������U��j�h�"d�    P���  V�  3�P�E�d�    ������\��������Pj�E�    ��B ��8�Q�B<��������Ѕ�u�����QP�B ����8�B�P�M�Q�ҡ�8�H�Aj j��U�h\$R�Ћ�8�Q�J�E�P�E��ы�8�B�Pj j��M�hP$Q�ҡ�8�H�A�U�R�E��Ћ�8�Q�Jj j��E�hH$P�ы�8�B�P�M�Q�E��ҡ�8�H�A��@j j��U�h<$R�Ћ�8�Q�J�E�P�E��ы�8�Bj j�h,$�M��PQ�ҡ�8�H�A�U�R�E��Ћ�8�Q�Jj j��E�h$$P�ы�8�B�H��(��e�V�E��ы�8�B�P�����VQ�ҍ�������P�K�������8P�B�M�Q�H����e�V�E��ы�8�B�P��`���VQ�ҍ�������P��������8P�B�M�Q�H����e�V�E��ы�8�B�P��P���VQ�ҍ�������P��������8P�B�M�Q�H����e�V�E�	�ы�8�B�P��@���VQ�ҍ�������P�s�������8P�B�M�Q�H����e�V�E�
�ы�8�B�P��0���VQ�ҍ� �����P�+�������8P�B�M�Q�H����e�V�E��ы�8�B�P�� ���VQ�ҍ� �����P����������M�Qh'  �E��� ��P��@���R�����VP��`���P�E��������P��p���Q�E��������P������R�E�������P������P�E�������P�����Q�E�������P�U�R�E��y�����P��0���P�E��e�����P������Q�E��Q�����P��P���R�E��=�����P��p���P�E��)�����P������Q�E�����P�E��> ��8�B�P������Q�E��ҡ�8�H�A��p���R�E��Ћ�8�Q�J��P���P�E��ы�8�B�P������Q�E��ҡ�8�H�A��0���R�E��Ћ�8�Q�J�E�P�E��ы�8�B�P�����Q�E��ҡ�8�H�A������R�E��Ћ�8�Q�J������P�E����E���8�B�P��p���Q�ҡ�8�H�A��`���R�E��Ћ�8�Q�J��@���P�E��ы�8�B�P�� �����@Q�E��ҡ�8�H�A�� ���R�E�
�Ћ�8�Q�J������P�E�	�ы�8�B�P������Q�E��ҡ�8�H�A������R�E��Ћ�8�Q�J������P�E��ы�8�B�P�M�Q�E��ҡ�8�H�A�U�R�E��Ћ�8�Q�E��E��JP�ы�8�B�P�M�Q�E��ҡ�8�H�A�U�R�E��Ћ�8�Q�J�E�P�E� �у�0������E����������   �M�d�    Y^��]� �U��E�MVW�   �;u��������s��th��8+�uE��������tQ��8+�u.��������t:��8+�u��������t#�� +�t�Ҹ   ���3Ʌ���_^��]�3�3Ʌ���_^��]���t$�m �����U��V���t$�m �Et	V�3 ����^]� ���������U����M�� ��A�@�X�A�@�X]� ������������U��E�@� �@����������������]��m ������������U�������E��������D�E{�ًM���������A���X�I�X]����P�P�]��������������U��M�U��"�E��A�b�X�A�b�X]���������������P�P��P(�P �P�P@�P8�P0�PX�PP�PH����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX��������U������P�M�P��P(�P �P�P@�P8�P0�PX�PP�XH���Q�P�Q�P�Q�P�Q�P�I�H�M��P�Q�P�Q�P �Q�P$�Q�P(�I�H,�M��P0�Q�P4�Q�P8�Q�P<�Q�P@�I�HD�M��PH�Q�PL�Q�PP�Q�PT�Q�PX�I�H\]� �����������U��M�U�A�
�E��B�I0���B�IH����A �
�A�A8�J���AP�J���X�A(�
�A�A@�J���AX�J���X�A�J�B �I0���B(�IH���X�A8�J �A �J���AP�J(���X �A@�J �A(�J���AX�J(���X(�A�J0�A0�J8���AH�J@���X0�A8�J8�A �J0���AP�J@���X8�A@�J8�A(�J0���AX�J@���X@�A�JH�BP�I0���BX�IH���XH�BP�I8�BH�I ���AP�JX���XP�A@�JP�BH�I(���AX�JX���XX]�������P�P��P(�P �P�P@�P8�P0�PX�PP�XH���������U��j�h�"d�    P��VW�  3�P�E�d�    �U�E�    ��8�H�I(R�E�P�ы���8�B�u�HV�E�   �ы�8�B�HVW�ы�8�B�P�M�Q�E�   �E� �҃��ƋM�d�    Y_^��]����������������U��UV���    �F    ��8���   �ARV�Ѓ���^]� ��������������U��UV���    �F    ��8���   �A(RV�Ѓ���^]� ��������������U��UV���    �F    ��8���   �E�I\RPV�у���^]� ���������̡�8���   �Q��Y���������������U���8���   �RD]��������������U���8���   �Rh]�������������̡�8�P@�B,Q�Ѓ����������������U���8���   �R|]������������������P�P��P(�P �X��$�@0    ����������X�X��$�������X���X �X(�������U��y0 ts��U�����Au���A�Z����Au�B�Y�A�Z����Au�B�Y�A�����z��Y�A �Z����z�B�Y �A(�Z����zZ�B�Y(]� �E��Q�P�Q�P�Q �P�Q$�P�Q(�@�A,�Q�A��Q �A�A$�Q�Q(�A�A,�Q�A�A0   ]� U��y0 �Et-�A��A �A�A(�A��$����������X���X]� ���P�P�]� ���������U��j�h1#d�    P��VW�  3�P�E�d�    �EP�M��E�    �� ���E�   � ��8�Q�u���BV�Ћ�8�Q�Bj j�WV�Ѓ��M��E�   �E� �� �ƋM�d�    Y_^��]��������U���V�u���O �]����e �]����{ �E��E�^�E��X�X��]������U��E� �@�@�E�E����������X���X]���������U���xV�uj ���! �@j�]Ћ��! �@j�]؋��! �@j �]����! �@j�]����q! �@j�]����b! �@j �]ȋ��S! � j�]����E! � j�]����7! � j �]����)! �@j�]���! �@j�]����! �@�E�u�E�E���P�ɍM�Q�]��U��E�R�ɍE�P���]����]��D�����^��]��������������U��V�u��u3�^]á�8���   �B(���Ѕ�t6���$    ���8���   �B(���Ћ�8���   ���B(���Ѕ�uԋ�^]����������������V����t}��8���   �B4���Ѕ�ui��8���   �B(���Ѕ�uR��8���   �B0���Ћ���t7�I ��8���   �B(���Ѕ�u;�t��8���   �B0���Ћ���u�3�^���������V����t}��8���   �B4���Ѕ�ui��8���   �B(���Ѕ�uR��8���   �B0���Ћ���t7�I ��8���   �B(���Ѕ�u;�t��8���   �B0���Ћ���u�3�^���������U���8�H@�U�A,VR�Ћ�8�Q�����B4j h�  ���Ћ�8�Q�B4jh�  ���Ћ�8�Q�B4jh�  ���Ћ�8�Q�B0jh�  ���Ћ�8�Q�B0jh�  ���Ћ�8�Q�B0jh�  ���Ћ�8�Q�B0jh�  ���Ћ�8�Q�B0jh�  ���Ћ�8�Q�B0jh�  ���Ћ�8�Q�B0j h�  ���Ћ�8�Q�B0jh�  ���Ћ�8�Q�B0jh�  ���Ћ�8�Q�B0j h�  ���Ћ�8�Q�B0j h�  ������$��8�Q�B,���$h�  ���Ћ�8�Q�B4jh�  ���и   ^]� ��U���8�H@�U�A,VWR�Ћu��j �΋��L �8�  j u��8�Q���   h�  ����_^]� ���L �8�  j u(��8�Q���   h�  ���Ѓ����_��^]� ���QL �8�  u*��8�Q���   j h�  ���Ѓ����_��^]� _�   ^]� ����U����  3ŉE���$��$��$�M��$VW�}�E��$�U��$�M�3Ʌ��E��U�~/�u�E�+����$    �T�ҍD�t���t:�u��;�|�_�   ^�M�3���^ ��]� �M�_3�3�^��^ ��]� �������U���,�  3ŉE���tXW��: ����uK�E�PW�; W��: ����t!��8���   ��4  j$�E�Phk� ���Ҹ   �M�3��b^ ��]ËM�3�3��R^ ��]�����U�����tW��8���   ��8  �U�R�U�Rhk� �Ѕ�t2�}�$u,�M�Q�U�R��7 ��P��H�V�P�N���V�Ƌ�]á`/�d/�h/��l/�N�V�F�Ƌ�]���������U����   ��8�HH���   SV�uj h�  V�҉E���8�HH���   h�  V3��҃���~K�u������F��U�'h�  R���^����F��g�^��F��g�^��8�HH���   �Ѓ�;�|��u��8�QH�B$���ЍM�WQ���AY P��<���SR������8�QH��P�B(����^[��]����������U���4�  3ŉE��E�U�E܋E�U��U�E�U�裏 ��u�M�3��\ ��]Ë�8���   SV�ȋBXW�Ћ؅�tY��I �ˍu��&�����M�P�U��H�M�P�E�P�U��8 ����t�M�Q�U�R���������u"3��������؅�u�_^3�[�M�3��\ ��]ËM�_^��3�[�\ ��]�������U���4�  3ŉE��E�USV�E܋E�U��UW�E�U��0t �؅�tr�u���t��8���   �B����;�uE�ˍu��R�����M�P�U��H�M�P�E�P�U���7 ����t�M�Q�U�R���������u"3����N����؅�u�_^3�[�M�3��C[ ��]ËM�_^��3�[�0[ ��]���U��j�h[#d�    P��   SVW�  3�P�E�d�    �} ��  �u�N��u3���F+����};��  �o  �ɋ]t�F+���;�r��^ �F�<� tS���-l  � �M�d�    Y_^[��]�k�p��  �}u�p ���u��h  �� ���E�������   �KhQ��t���R���������8���   P�B|���E�    �Ћ�8�Q�J��t���P�E������у��{�?�����8���   �u��P����=�����   �Ej P��葵 ��   �}��KHQ��l���R�������M��P�U��H�M��P�U��H�M��P���ˉU��: �؋���؉E��E��: �U�M���Q�M�R�E��?� ���1  3��M�d�    Y_^[��]Ë��L: �؋���؃�P�� ���4: �؋���؃�P��� ���U܍E��U�P���]��� �KHQ��T���R������M̋P�UЋH�MԋP�U؋H�M܋P���E�P�ΉU��L� �} u<�M�nj  ��u0j h�  ���|� �����;����KQ�M�j  �R���l� �W����9 ��|L���9 �M����  ;�}7j h�  ���,� ������������9 �MP��i  � P���� ��u��MQ�M�i  ��S�0�]��)4 ������   �E���  3ۅɉM�~.���  ���I �U�RW�f�������u����p;]�|�E�M�;��_����}$�M �UWQ�MR�USQRP�EP�w����؃� ��tf��8���   �B����=���u'�Mj SV�h� ��聲 �ƋM�d�    Y_^[��]Ë�8���   �B4����j P�������PS�i�}$��8���   �B����=���u$�MV�� �������ƋM�d�    Y_^[��]Å�t��8���   �B4����P�]������3�j PW�MV�	p �ƋM�d�    Y_^[��]������U��QSV��W���7 ��tb�FP�E��2 ����uX�E���  3���~(���  ����E�PW���������u
����p;�|�E;�}k�p��  ���>7 ��u�_^3�[��]�_^�   [��]������U��j�h�#d�    P��h�  3ŉE�SVWP�E�d�    �E�M�U�}��P  �EЋE�MԋM�U؋U �E܋E$�M��M(�U��U8�E��E<3ۅ��M��U��E�~5��L  �Eă��EȋUȍM�QR��������u0��   E�Eȃ�;�|�3��M�d�    Y_^[�M�3��UU ��]ËE����tp��8���   �P4�ҋ؅�tY��$    �ˍu��������P�M��H�U�P�EЉM�P�M�Q�U�����������   ��8���   �P(���ҋ؅�u��u�3��ẺE��F3�;���  �]��I �FE�9�`  ��P�M��H�U�P�M�U�]���  �]���\  u��E��^P�KQ����������8  ���Fb ���)  �}4 t5�V�Nh�  ���ĉ�V�H�N�P�H�M��/������	������3��U��E,�M�R�U�Q�M�P�E����$R�U�PQRWV�X  ��,���E���   �M̅�u,��8���   �ȋB��=  t�MȉM��   �M̅�t1��8���   �P��=  u��8���   �E̋MȋRDP���Qh  �� ������u�E�P�� ���0�M̅�t��8���   �PDV�ҡ�8���   �MȋBDV�ЉűE��E��   ��;�`  �E�������u�3ۋE��E���;F�E��>����N(Q�U�R�a�������8���   �M�P�B|�]��Ћ�8�Q�J�E�P�E������э~�ũ�������u�9unh  ��� ��;Éu�U�R��� ��������8���   �M��RDQ����h'  �S ��8���   ���P�B|�Ћj�� �j芾 ��8���   ��M̋RDP�ҋE����������������U��j�h�$d�    P���  SVW�  3�P�E�d�    �ك}�}�5  ��8�H�A�U�R3��Ћ�8�Q�J�E�P�u��эUR�E�P�M�QV�E���) ����t#����} u�UR�E�P�M�QV��) ����u�j ����= ��8�8�  �B��  �P�M�Q�ҡ�8�H�Aj j��U�h&R�Ћ�8�Q�J��d���P�E��ы�8�B�Pj j���d���h&Q�ҍE�P��d���Q��8���R�E�������M�QP��(���R�E��������@P��H����E��C� ��h�%�������E��� ��������P�E��ۛ WP�����Q�E��� VP��H���R�E�	�׋ ��������E��e� �������E��V� �������E��G� ��H����E��8� ��8�H�A��(���R�E��Ћ�8�Q�J��8���P�E��ы�8�B�P��d���Q�E��ҡ�8�H�A�U�R�E��Ѓ�行 �Eh1D4ChCD4Cjjj��H���Q��Ȉ]�軌 ��j h�%��   �M�����j h�%�M��E��q����U�R��H����E��.� P�E�P��t���Q�E��i����U�RP�E�P�E��W���P�E��� ��8�Q�J�E�P�E��ы�8�B�P��t���Q�E��ҡ�8�H�A�U�R�E��Ћ�8�Q�J�E�P�E��ы�8�B�P�M�Q�]��҃�0�}  �M�����j h�%�M��E�����h�%��,����E��ׅ ��h�%��d����E���� ��������P�E�诙 WP������Q�E�轉 VP������R�E�諉 ���M�Q���E���� P�U�R��t���P�E� �4����M�QP�U�R�E�!�"���P�E�"� ��8�H�A�U�R�E�!�Ћ�8�Q�J��t���P�E� ���E���8�B�P�M�Q�҃�(�������E�貅 �������E�装 �������E�蔅 ��d����E�腅 ��,����E��v� ��8�H�A�U�R�E��Ћ�8�Q�J�E�P�]��у��UR�E��� ����H����E    �E��#� ��8�H�A�U�R�E� �Ћ�8�Q�J�E�P�E������у��   �M�d�    Y_^[��]� �P�M�Q�E� �ҡ�8�H�A�U�R�E������Ѓ��M�UWQR���3 �M�d�    Y_^[��]� �������������U��j�h�$d�    P���   SVW�  3�P�E�d�    �]����$3����u����E��$�ʉu�ݝp����u��ɉu�ݝx����]���$�������]����]��]��u��E�%�uЉuԉu؋���   �M�Q�U�R���E��Ѕ���  �����詹 �����   V��������$P���E��҅��u  ��Px���҉E�3Ƀ��   ����h&h�  hD����Q�m ����P|��V�ωu��E��҅��  �E�P�M�Q����� ����   3�9M܉M���   �E��E����U��D�������A��   ����������   ������z�����U���������z������3�8U���;�U�i�����Eݝh�����ݝ`������I �E��Eă���H�����ܵh���܍`������$P�( P�M��k  ��;�u�~��E��M��E��u��E� ��u������E� �������؃�;M܉M��������؅�t	V�� ��3�������E��}� �}���   ����   ���Ѕ��}�t���;���   �u���E��H����F�Q�F��p����������������ݝH���ݝP���ݝX������������u�3�9u�t3�E��}܅p����E�܅x����E��E���$����������_�_���E�P���P�9u��E� �E�%t�E�;�tVP�M��%�uЉu؉u�9u��E������E��$t�E�;�tVP�M���$�ǋM�d�    Y_^[��]����������������U��j�h%d�    P��   SVW�  3�P�E�d�    �ً}3�;���  ;�t�]��VV��� ���E���;��k  ��8�HH���   h�  S�҃���u=��8�H@�Q,S�ҋ�����   �����ҋ�8�Q�����P�B0h�  ����3��E��$�uԉu؉u܉u��E�%�uĉuȉű���   �E�P�M�Q���E��҅���  ��h����ε �����   V����h����$Q���E��҅��l  ��Px���҉E�3Ƀ��   ����h&h�  hD����Q� ����P|��V�ωu��E��҅��  �E�P�M�Q����� ����   3�9M�M���   �E��E����U��D�������A��   ����������   ������z�����U���������z������3�8U���;u�U�\�����E�]����]���E��E����P������u��M����$P�]	 P�M��Dg  ��;u�u�~��E��M��E��]��u��E� ��]��ۋu����E� �������؃�;M�M��$������؅�t	V�� ��3���h����E��� 9u�/�M��E� �]  �M��E������ 3��M�d�    Y_^[��]Ë�8�QH���   h(  S�Ћ�8�QH�E싂�   h�  S�Ћ�E䋂�   �����Ѕ�t�u؃���u���M؉M��E�U��P�E�P���e� ��8�QH���   j h�  S���E��3ۃ���   �U�����3ɍR���Ѝ�    �}��9��`�D9���`���D9����������������Z����Z��Z��}��D9��D9��D9����������������Z����Z��Zȋ}��D9��D9��D9����������������Z����Z��Z��}��D9��D9��D9����������������Z����Z��Z��R����}�u�;�}J�U�Ӎ[ɍRɍЋ��+Ӌ]�����D������D����������������X����X��X�uΡ�8�؋HH�U����   j h(  R�ЋM�؉t������   �����ЋM�����؉D��3�9u��E� �E�%t�E�;�tVP�M��%�uĉủu�9u��E������E��$t�E�;�tVP�M���$�E��M�d�    Y_^[��]������U��j�h�%d�    P��t  SVW�  3�P�E�d�    3��}��E�%�}̉}Љ}ԋ]�K��P(�}��҃��u�1  ��  ���r  ��t���7  �E0� �,  �CP�� �������  ��8�Q���   jh�  ���Ѕ���   ��8�Q���   j h�  ���Ћ�8�Q���   jh�  �����E �����$PW3������؃��ۉ]���   ��8�Q���   jh�  ���Ѕ�tu��8�E �Q���   ���$jh�  ���Ѓ�P��d���Q�������݅l����ȃ�݅d�������݅t��������C ��&����AuS��d����;���������  �EЅ���  3�3�3�;��M�M�}��M�M��}  �  �SR�
� ����;�t�h  ��� �؃��ۉ]�t��E ���$����8���VP�������8�QH��P�B�����q�����8�Q���   jh�  ���Ѕ��W����KQ�� �����C����U�Rj����l ���.����E,� �#����� ��  =   �  =   @t�E0� ������CP�q ��;ǉE������3�ǅl���,%��p�����t�����x���h�  �E��ڿ �؃�;߉]�u��l����E� ��Y  ������&���$jj���S� ���,�����8�Q���B4jh�  �����E �]���K�$Q�U�R�����E ���C �$P�M�Q�t����E��e���8�E����e��������E�Q�e�h�  �ʋ�ݝ����ݝ����ݝ�����B�PH�ҋ�� ����   �$�h\ ��8�P�B0j h�  ����j h�  �o��8�Q�B0jh�  ���Ћ�8�Q�B0j h�  �����8j ��8�Q�B0h�  ���Ћ�8�Q�B0jh�  �����j�΅�tjh�  ��8�Q�B0���С�8�8�>  |�P�B0jh�  ���Ѝ�l���Q���� ����  ��8�B���   jh�  �������U����U��E��]��g ����   ��8�P���   jh�  ���Ћ�8�Q���   jh�  �����E 3�9�t����������$P��#�p����	Q3�������8���؋B���   jh�  �����E 3�9�t����������$P��P���P��#�p����	�����  j j �4� 3���9�t�������   ���8�Q���   jh�  ���Ћ�8�Q���   jh�  �����E ���$��PW��l����P  �Q���������}� tM��8�B���   jh�  �����E ���$��PW��l����O  ��h���Q��������P�M�������;�t����D����}� t8�M��� �E��E����U��$R�� ���P������ ���]��@�]��@�]��������+������������ �����Q�M���$�	 ��tG����������$R������P�*���������Q������R��@���P�����   ������������8�QH�B$���Ѝ�����QP������R�������8�QH��P�B(���Ѓ}� t1�E����E������E������= ��&����AuS�}��R�������t�M�Q��������l����E� �aU  �]�������SR��� �����������h  ��� �؃��ۉ]�������E ���G�$P������Q� �����8�RH��P�B(�����E �M0�U,3�9E(Q�MR�U��P�E���$VQ�MR�WPQ�G���̉�P�Q�P�@�Q�A��������8���8������������8�QV�ȋBph�  ��������8�Q���   jh�  ���Ѕ�������KQ��- �����E�������U�R�M��\  ������d$ 3ɋE̋4��V�F U�E�;�u���A[ ��u3���   �}� u���G[ ���E�    t�E�   �}� u���H[ ���E�    t�E�   ��;]�|��}��u(3�3�;��u؉}���|�����X�����\�����`�����   �M�U�QR���ߩ ��u;�}� �E������E�%t�E̅�tj P�M��$%3��M�d�    Y_^[��]á�8�HH���   j hO  V�ҋ���8�HH���   j h'  V�}��ҋ؃���|�����E�M�PQ�!� �������u��f����}� t?��u;�U�WRhO  ���f� ���E�u#�M��E�������Q  3��M�d�    Y_^[��]Ã}� t��u�E�SPh'  ���!� ����|���t��}� ��  �]�j Sh2  ����� j S��h2  �Ή�`����� �M�j Q��h2  �Ή�\����ʦ ������X����[������S������K���j h�&�M�苽����8���   �Px���E��ҍM�QP�U�R������P���E��7�����8�H�A�U�R�E��Ћ�8�Q�J�E�P�E� �у�j h�&�M�������8���   �Px���E��ҍM�QP�U�R������P���E��������8�H�A�U�R�E��Ћ�8�Q�J�E�P�E� �у�j h�&�M�詼����8���   �Px��Έ]��ҍM�QP�U�R������P���E��T�����8�H�A�U�R�]��Ћ�8�Q�J�E�P�E� �у��������<�����8�BH�}؋��   3�Sh�  W�]��у�9]ЉE��]���  �E��Ű<�3�9G�E�~`�u��[�u�E��4����    �GE��U�� R�@�������@�E ����������^�^� ����E�E��E�����;G�E�|���8�HH�U؋��   j h�  R�Ѓ��  �E��E�    ~n�u����E�    ��OM�M��,/ �U��J˄���Rt�Ӊ�N�F�ӉUċU��R�Ӊ�UĉV�N�E��F�E����;G �E�|��}� �\  ���V ���M  �M��z� ��������  �E�    �,  �M��x&�u������T2�I�U�t��U�B��O,+Í@�����@�@������A ��f�F���A ��f�F���A �U�f��B��O,+Í@�����@�@�����A ��f�F�A ��f�F�A �U�f�F��O,+Í@�����@�@�����gA ��f�F�\A ��f�F
�QA �U�f�F�B�O,+Í@�����@�@�����*A ��f�F�A ��f�F�A �E�f�F�E����E���;G ������؋�|������r  ���@U ���c  ���ݕ���ݕ ���ݕ����ݕ ���ݕ���ݕ���ݕ8���ݕ0���ݕ(���ݕP���ݕH���ݝ@���臞 ���E������  �E�    ��   �U�E����t���   �N�+ˋȋL��M��N��U��E�ݝ����+��E�ݝ �����ݕ����ȋL��M���U��E�ݝ���+��E�ݝ���ݕ ����ȋL��U��E�ݝ(����M��E��Nݝ0���+�ݕ8����ȋD���8�U��E�ݝ@����E��E�������ݝH���P�E�ݝP����QD�M��R0�Q�M�Q�ҋE�������;G �E���������S ����   ��X����[� ��\����E��M� ��`����E��?� � �E�    �o   �MċU�+�+��4��UĉE��	��$    ����  �M����M��� �]��M��!� �]��M��6� �E��UċE��2�E����^��\0��E���;G�E�|��E��O _M��;EЉE��:����}؋�8�B�M���   jh�  �҅���   �M����? ����   �E�P�����������M�Q������R�. ��8�QH��P�B(���Ћ�8�QH���   h�  W3��Ѓ���~G�u������F�h�  �e�W�����^��F��e��^��F��e��^��8�QH���   �Ѓ�;�|���8�Q�]���   3�Vh�  ���Ѕ���   �u��u��u��u��u��M��E��u��}��� �p&��8�Q���   ���$h�  ���E�	�Ћ�8�Q�B,���$h  �M��Ћ�8�Q�B0jh  �M��Ћ�8�Q�B0Vh  �M��Ћ�8�Q�B0Vh  �M��ЍU�R�M�h�   �M�� ���M��E���� �M��E� � �h&���$Vj���;� ��8���   �BVj���Ћ�8���   �BT���Ѕ�u�}܃}� tO�}�O Q�U�R��������8���   �u�P�B|���E�
�Ћ�8�Q�J�E�P�E� �у��������}� �E������E�%t�E̅�tj P�M��$%�E܋M�d�    Y_^[��]ÍI 8L WL �L �L ��������U��j�h�%d�    P�� V�  3�P�E�d�    h'  �@�  ���8�H�A�U�R�Ћ�8�Q�J�E�PV�ы�8�B�P�M�Q�E�    �ҡ�8�H�Aj j��U�h�&R��j �M�Qh�� h   �U�RhS� �E���� ���8�H�A�U�R�E� �Ћ�8�Q�J�Eԃ�@P�E������у��ƋM�d�    Y^��]��������������U��j�h�%d�    P��SV�  3�P�E�d�    �u3�;��9  ���] ��8���   �BSh  @j�����E�   �]܉]��]��]�]�Ή]��F �؅�tV��I ��8�Q@�BS�Ѓ��u"�E�����|jjjP�M��2I  ��t�M�����8���   �P(���ҋ؅�u�3�9]�~t��3�这  ��v4�O��t�G+���;�r�1 �G���U�;�t�σ�苙  ;�r̋�耙  ;�s �E���Q�Mj-�K\ �U���P�o� ����;]�|��M�\ �}� �E�����t�M�Q�6�  ��3��M�d�    Y^[��]�U��j�h
&d�    P��$SVW�  3�P�E�d�    �u3�;�u3��M�d�    Y_^[��]Ë��t[ ���-E ;ǉE���  �u��3�趘  ��v3���N;�t�F+���;�r�0 �F�M�9�t�΃�胘  ;�rϋ��x�  ;��  �E�   �}Љ}ԉ}�}܉}؋M�}��D ��3�;��}���  ��}�9}��\  ���+�  ��v8��$    �N��t�F+���;�r�"0 �V�E�9�t�΃���  ;�rϋ���  ;��
  �M�W�G� ����   ��8���   �Bx���Ћ�8���   �M��؋Bx�Ћ�8�Q�ȋBxS�Ѕ���   �E����|jjjP�M��F  ��t�Mԉ<��M�C ���E����   ��8�BH���   3�Wh�  S�ы�����tGj ���ʏ ;E�u�MVj*��Y �U�R���Ϗ ��8�HH���   ��Wh�  S�ҋ�����u��}�������؅�u��u�}��8���   �B(����3�;ÉE��y���3�9]�~(�Mԋ��MRj-�Y �Eԍ�Q�� ����;u�|�9]��E�����t�U�R�s�  ���]Љ]ԉ]�]܉]�3���8���   �M��B(��;ǉE������u����X �   �M�d�    Y_^[��]�U��j�h�+d�    P�DL  ��6 �  3ŉE�SVWP�E�d�    �E�M�U�� ����E������������C:  ����x���t
j ��  ����ȸ�����	 �������(���P�E�    �?b ��8�Q�Bdj ��(����E���h&��h)  �{hD�W�K�  ��8�Q��j ���BhWV��(�����h�'V��ȸ��� ���	 ����t	V��  ����u6��8�Q�J��(���P�E� �у���ȸ���E��������	 ����]9  Wj�������	 �������E��sH j �����R�������E��kf W�����	 ����uT�������E��J ������E��	 ��8�H�A��(���R�]��Ѓ���ȸ���E������b�	 �������8  ��x��� �   t	S��  ��j ��������� ��u9�������E��AJ ������E��B	 ��8�Q�J��(���P�E� ��뀋E�ȃ� ǅԸ��    ��l�����   ���   �������? ����и����   ���    ��и���ύ�����������U��H�M�P�U�@�M�Q�E�� ����t-�U��M�j ���ĉ�U�H�M�P�H��x����-� ��u��и��3����������и��u��%��t!h'  ���  P�, ����t
ǅԸ��   ��8�B@�� ����P,Q�����8ݝ�����Q��j ��ظ���ȋ��   h�  �Ѕ��  �� �ȉ������(���������E���   �$��� ��'j��   j��   j��   j�   j�   ��'j�   j�   ��'j�   ��'j�   j�   ��'j�x��'j�n��'j
�d��'j
�Zj
�Tj	�Pj�Lj�H��'j
�@�x'j
�6�p'j�,�h'j�"�`'j��X'j�݅0���j�j ����$��~ ��l��� tl��8�Q@������B,W�Ѓ�h��hE  ��輺 �������Q���l ����   �����VR�G� ݝ�����������R�E��� ��   �����Ph����������������8�Q@������B,W�E��Ћ�8�Q��V�ȋ��   hE  �Ћ�8���   �
������P�E��у������R�E��M �w��ظ��h��hE  �� Ph��������腼�����8�H@������Q,W�E��ҋ�8�Q��V�ȋ��   hE  �Ћ�8���   �
������P�E���3���9�Ը����������   h  �#� �������������40  �������д��P�] ��д���E��_^ ������Q��д����] ��8���   P�B|���E��Ћ�8�Q�J������P�E��у�j j j V���< ��д���E��l[ 3���8�B��ظ�����   jh�  ��9�Ը������и���{  ��8�P��ظ�����   jh�  �Ѕ��V  9�P���������D  ������	��$    ����L���������<�<� �����|  ��X  P������Q��������8���   P�B|���E�	�Ћ�8�Q�J������P�E��у�������R��0���P����  ����Z � �@������@Q�ʋ�ݝ���ݝ���ݝ����R  � ��̶���@R�@����ݝ����ݝ����ݝ������� � ���@�@��������PݝH���ݝP���ݝX����� � ������@Q�@������݅����R�ˍ�H�����P�ɍ�ȷ����ݝȷ��ݝз��ݝط��Q�������?�����8�RHP�B0���Ѝ�p���Q���B ��p����u_ ����   ݅��������p����$R�����P莼��݅������P���������$Q����� P��H���R�c�����P��ȷ��P����P荴��ݝ������ǅ���   h�  �������E�
�� j �����QP���E��q �������E�
�� ��8���   ������Q�E��҃����m� ��tK�E�   �E�   h�  ��|����E��W j �M�QP���E�� ��|����E��V �M��5  ǅ@���   ǅH���    h�  ��X����E�� j ��@���QP���E��~ ��X����E�� ��8���   ���@���Q�E��҃���`���P��� ݅`����   ݝ����������h�  �������E�� j ������QP���E��6~ �������E��
 ��8���   �������Q�E����P'ݝh�������`���h�  �������E��# j ��`���QP���E���} �������E��
 ��`�����8���   �Q�E��ҋ������������j j PV�8 ����������(  ��;�P���������������и��3������������������9�Ը���]���
  ���y	  9������������
  ������Ƹ ��3�;���  ������������<�OQ������R諸������8���   P�B|���E��Ћ�8�Q�J������P�]��у�ǅ���   ǅ����   hn  �������E��� j �����RP���E��x| �������E��� ��8���   ������R�]��Ѓ��E�   �E�   h�  ��|����E��k j �M�QP���E��| ��|����E��j ��8���   ��M�Q�]��ҍG(P��p���Q�C�����P��8����Ĵ���� ���h4  ��X����E��� �� ���j RP���E��{ ��X����E��� ��8���   ���8���R�]��Ѓ�j�jj ��蝲 ���?  i�X  Gh�x! �,  �H�� ����� ���  h�  �B �����������   h�  ��h����Q �� ���Q��Զ��R�E�躶����P�������E���S P������E����������j P��h���P�E��z ��8���   �
�����P�E��у��������E���S ��8�B�P��Զ��Q�E��҃���h����]��� ��8���   ��������   j P���ҋ��R�����8�Q������RpQh@  ������'�_P����A��   ǅ@���   ǅH���    h�  ��`����E� �* j ��@���QP���E�!��y ��`����E� �& ��8���   ���@���Q�]��҃�ǅ����   ǅ����    h�  �������E�"�� j ������QP���E�#�ly �������E�"� �������  �O0��� ��8���� 3�;���ǅ`���   ����h����$h�  ��p����]��P j ��`���RP���E�%��x ��p����]��M ��8���   ���`����   R�]��ЍG0P��p���Q������P������蠱���� ���h  �� ����E�&�� �� ���j RP���E�'�x �� ����E�&�� ��8���   �������R�]��Ѓ�ǅ\���   ǅd���   h�  ��8����E�(�n �E�)j ��\���QP���x ��8����E�(�j ��8���   ���\���Q�]��҃�ǅ����   ǅ����    h�  ��P����E�*� j ������QP���E�+�w ��P����E�*� ��8���   �������Q�]�����ݝD�����ǅ<���   h�  ������E�,� j ��<���QP���E�-�Iw ������E�,� ��8���   ���<���Q�]��҃�踉 �P�����H'��% �@'ǅ���   �8'ݝ����E�.h�  ��$���� j �����QP���E�/��v ��$����E�.� �������8���   �Q�]�����'�_X��������  ǅ���   ǅ$���   h�  ������E�0� j �����QP���E�1�Dv ������E�0� ��8���   ������Q�]��ҍG8P��p���Q�k�����P��|��������� ���h`	  ������E�2�" �� ���j RP���E�3��u ������E�2� ��8���   ���|���R�]����GXݝ4�����ǅ,���   ha	  ������E�4� j ��,���QP���E�5�fu ������E�4� ��8���   �]����,���Q���G@ݝT�����ǅL���   h�  �������E�6�S j ��L���QP���E�7��t �������E�6�O ��L����Rǅl���   ǅt���    h�  ������E�8�� j ��l���QP���E�9�t ������E�8��  ��l�����8���   �Q�]��ҋ������j ���?. P�9�����PV���. �� ���P������� ����%C  �����������   ��;���������������  �����;�t	P��  ��������������������������E��7 ������E��� ��8�Q�J��(���P�E� ���!  ���E  9�����������3  ������D� �����#!  ������������<�OhQ������R�+�������8���   P�B|���E�:�Ћ�8�Q�J������P�]��у�H��p���WR舯����P��8����	�����h4  ������E�;�C j WP���E�<��r ������E�;�E�  ��8���   ���8���R�]��Ћ������j ���, P脰����PV���- �� ���Q������� ����pA  ����������p��;���������������3��������� ���PQ�������� ����<  ��8�B��ظ�����   j�=h�  �ψ]���9�Ը���������  ;���   3�9�������   3ۃ�����������T�Du+j����̉�P�Q�P�@�Q�A������������'���̉�P�Q�P�@�Q�A���������������t'��������t������+���;�r�� �������4�����p;������X���3�3ɉ��������������9�Ը���E�m��   ��8�B��ظ�����   jh�  �҅���   9������������   3ۍ�    hF  �f� ��3���;��� ����D  �������<�OQ������R�x�������8���   P�B|���E�n�Ћ�8�Q�J������P�E�m�у���������� ���R��ܸ���?  ��������� ;�����������Y���3������9�x���tj���  �������9� ���������������,���ǅl���   ������f  �� �����I �����������^�ˉ�t���� ���   ��8�B��ظ�����   j h�  �҅�t2��� ����  �C k�p�����������Q�!���������  ��Ը�� ��  �V�Nh�  ���ĉ�V�H�N�P�H��葴�����X  ��8�Q���   jh�  ���Ѕ������9�����������������T�����������T���h�  �4�f� 3���;ǉ�����  ���ݕȷ��ݕз��ݝط���H� �H��   ;��6
  �$� � ǅ|���   ǅ����   h�_ ������E�>� W��|���Q�����P�E�?�an ������E�>��  ��8���   ���|���Q�]�����	  ǅ$���   ��,���h�_ �������E�@�O W��$���Q�����P�E�A��m �������E�@�H�  ��8���   ���$���Q�]����c	  ǅ\���   ǅd���   h�_ ������E�B�� W��\���Q�����P�E�C�m ������E�B���  ��8���   ���\���Q�]��҃����o ���   �����ݝ����h�_ ������E�D�o j �����Q�����P�E�E�m ������E�D�g�  ��8���   ������Q�]���݅����Q��p����$P���up P��H���Q�h���P袡��ݝ������������h�_ ������E�F�� j �������E�GR�����P�l ������E�F���  ��8���   �������R�]��Ѓ�3���  ǅ����   ǅ����   h�_ ��$����E�H�l W������Q�����P�E�I�l ��$����E�H�e�  ��8���   �������Q�]���݅����Q�������$P���so P������Q�f���P蠠��ݝ������ǅ����   h�_ ������E�J�� �����W������RP�E�K�k ������E�J���  ��8���   �������R�]�����  ǅ����   �����h�_ ������E�L�p W������Q�����P�E�M�k ������E�L�i�  ��8���   �������Q�]����  ǅԵ��   ǅܵ��   h�_ �������E�N� W��Ե��Q�����P�E�O�j �������E�N���  ��8���   ���Ե��Q�]��҃����7l ���   �����ݝ���h�_ ��4����E�P� j �����Q�����P�E�Q�7j ��4����E�P��  ��8���   ������Q�]���݅����Q�������$P���m P�����Q艦��P�Þ��ݝ�����������h�_ �������E�R�  j �������E�SR�����P�i �������E�R���  ��8���   �������R�]��Ѓ�3��  ǅ<���   ��D���h�_ ��t����E�T� W��<���Q�����P�E�U�9i ��t����E�T��  ��8���   ���<���Q�]��҃�ǅ���   ǅ���   h�_ ��T����E�V�% W�����Q�����P�E�W��h ��T����E�V��  ��8���   ������Q�]����9  �   ��l�����t���h�_ ��4����E�X� j ��l���Q�����P�E�Y�ah ��4����E�X��  ��8���   ���l���Q�]��҃���ĵ��ǅ̵��   h�� ��$����E�Z�Q j ��ĵ��Q�����P�E�[��g ��$����E�Z�I�  ��8���   ���ĵ��Q�]���݅����Q��(����$P���j P�����Q�J���݅��������@����$R����i P��p���P�#���P�]�����$��ǅL���   ݝT���h�_ ������E�\� j ��L���Q�����P�E�]�7g ������E�\��  ��8���   ���L���Q�]���݅�����$����3�݅�����݅�������ݝȷ����ݝз��ݝط���m  �   ��|���������h�_ ��D����E�^��  j ��|���Q�����P�E�_�f ��D����E�^���  ��8���   ���|���Q�]��҃�������ǅ����   h�� �������E�`�  j ������Q�����P�E�a�)f �������E�`�z�  ��8���   �������Q�]���݅����Q��X����$P���Hh P�����Q�{���݅�������������$R���Qh P������P�T��������Q舚��ݕ������$���   ݝܶ����Զ��h�_ ��d����E�b��  �����j ��Զ��RP�E�c�[e ��d����E�b��  ��8���   ���Զ��R�]��Ѝ�����Q����ܵ�����������ݝ����h�_ ��h����E�d�>�  �����j �����RP�E�e��d ��h����E�d�6�  ��8���   ������R�]���݅����܅�����݅���3�܅����݅���܅������$��������ݝȷ��ݝз��ݝط��������Q��� ��9�����v  ������R����g � �@��݅��������ݝh�����ݝp����H������Pݝ �����g � �@�@݅��������ݕX�������ݕ|���������ݕ������݅p�������݅ ���������ݝ8�������݅h�����������ݝ����������������ݝ`����������������^ ����������D{4������݅h�����݅p�����݅ �������ݝH���ݝP���ݝX������ݕX���ݕP���ݝH���݅8�����݅��������݅`��������� ݅8�����݅������݅`���������������D{&������������������ݝ����ݝ����ݝ�������������ݕ����ݕ����ݝ����݅X�����݅|�������݅���������b ݅X�����݅|�����݅����������������D{&������������������ݝ���ݝ���ݝ������������ݕ���ݕ���ݝ���������Q���e � �@��H����@R݅������������P�ʍ������Q�ʍ�p���܅ȷ��R݅з����������݅ط����ݝp���ݝx���ݝ����躗����8�QH�����P�B(�Ћ��nd ݝ@���ǅ8���   hQ�  �������E�f��  j ��8���Q�����P�E�g�aa �������E�f��  ��8���   ���8���Q�]��҃��� ���P���'d �����ޫ ݝ�������� ݝ|������� ݅����ݝp���݅|���ݝx�����8ݝ����3���������������   �R��p���P�����Q�҃�h�_ ��H����E�h���  W�����Q�����P�E�i�` ��H����E�h���  ��8���   ������Q�]��҃����g ݝ����ǅ����   h�_ �M��E�j�v�  W������Q�����P�E�k�` �M��E�j�r�  ��8���   �������Q�]��҃����^a P������P衛������8���   �����P�B|�E�l�Ј]���8�Q�J������P�у�����` ��u�����P��m ��������и���������   WRPQ�����R�����������P������QR�s������� ��tR��8���   �B����=��������uj j WQ������ �����V��[ �+��8���   �PHV�������������j j WP�q �������T����  ��;����������������a���������;�t	P�W�  ����������������ĸ���r��������;�t	P�-�  ��������;ǉ��������������t	P��  �������;ǉ�������������ĸ��t	P���  ��������������������������E��! ������E��� ��8�H�A��(���R�E� ���  3�݅���������R��ظ�������QP���������$RWP��,���Q������RV�S�����,��������{  ����ݕ����������ݕ����P��ݝ�����Z� ��t������� ����  �$�D� ��8�Q��ظ�����   3�Sh�  �ЋO �����������k�p������������DH��T�����T���躧 ��T����]��̧ ��T���ݝH����ۧ ݅H����E�ݝ����ݝ����ݝ�����=  �wP��ǅ����   �g� �]���}� ݝH�����萧 �������   ���. �� t��t�O ������k�p�D0��G(��G ������k�p�D0������i��   �D(��<�����<���ǅ����   �� ��<����]���� ��<����f��8�Q��ظ�����   j h�  �ЋO �����������k�p������������DH��$�����$����z� ��$����]�茦 ��$���ݝH���蛦 ݅H����E�ݝ����ݝ����ݝ����3ۍ�����Q���@~ ����
 ���r
 ����
 ��tS�������   Sh�  ���]j ;��V  ��8�J@�Q,P�ҋ��8�P�B0��jh�  ����Sh�  �]Sh�  ���j ;���  ��8�Q@P�B,�Ћ�8�Q�����B0jh�  ���Ћ�8�Q�B4jh�  ����Sh�  ��8�Q�B4���Ћ������и����u\9������  Sh�  ���i ��3�;��i  �����;ʋw t������+���;�r��� �������Q���^` �  ����  ����	 ���7  �O(;��,  �����;�u3��������+���;��  Sh�  ����h ��;��P  �W(R������  � P����_ h�  ���������  ǅ����   ǅ����   S������Q������R���E�p�vY ��8���   �������R�E�o�Ѓ��������E�m��  h�  ��|����z�  �0'ݝ@���ǅ8���   S��8���Q��|���R���E�r�
Y ��8���   ���8���R�E�q�Ѓ���|����E�m�>�  �]  ��� ���N  ������A  �O ������k�p�\0���'  �������t������+���;��
  �����j h�  �g �����f  S������0  � P���^ h�  ��X�����  ǅ���   ǅ����   j �����Q��X���R���E�t�X ��8���   ������R�E�s�Ѓ���X����E�m�K�  h�  ��`�����  �0'ݝܶ��ǅԶ��   j ��Զ��Q��`���R���E�v�W ��8���   ���Զ��R�E�u�Ѓ���`����E�m���  3�ǅ�����$�����������������������;��E�w�T  �����+����C  ;������7  ������Q��t���� ���  3�9������  �����������������4�����   ��u3����+���;���   ��t��+���;�r�K� ������������    �< ��   ��t	+���;�r�� �������8��J@�Q,P�҃�h�f h�  ���&� ��j t�����Q���� �;h�&�������|��������R�E�x� �  ��8�H�A������R�E�w�Ѓ�������������;������������������и���������t���WQ�H RQ�����R�����������P������QR�ڛ����3ۃ� ;�t@��8���   �B���Ћ�8���   =����BHuW���������V���TR �V���8���   �BHW�������9������E�mǅ�����$t*������;�t SP��������$��������������������x��� tD���������t���ۅt���ڵ �����&� �   +�;�l���~Q��l�����  ��������� ��������   ;� ���������� �������������3�������3�9�Ը����  3������;���  ��+���;���  �ʋ���8�� ����J@�Q,P�҃�h�f h�  ���� ;��L  ���5� ���=  ��8���   �B4����WP�ԑ���� �����PSQ������} ��������`��������;�t	P��  ��������;É��������������t	P�Z�  �������;É�������������ĸ��t	P�5�  ��������������������  �����;�t	P��  ��������;É��������������t	P��  �������;É�������������ĸ��t	P���  �����������������������������;�tP藺  ��3ҋ�����;��������������tP�p�  ��3ҋ����;�������������ĸ��tP�I�  ��3҉����������������������ܸ���  �������  �������  �������E��� ������E���� ��8�B�P��(���Q�E� �҃���ȸ���E�����萲	 �������  ��ܸ���  �������  ������  ������� ���R�dr ����������D��������;ы�v�<� ����������;�v�'� �����;�t'+����ɍ�    �<0~PSPV�|� �������3�9�Ը��uA��8�P��ظ�����   jh�  �Ѕ�t �����V�����������QV�x�����3�9�x���t
jZ���  ����������� 9�x���t
jd��  ���E�  ��8�B�P�M�Q�҃������;ǳy�]���   P������P�����P������h'  Q�E�z��  ������8�B�P<�M��E�{�ҋ�8�Qj�j�VP�BL�M��Ћ�8�Q�J������P�E�z�ы�8�B�P������Q�]��҃�9�����&  ��8�P�B<�M��Ѕ���   ��8�Q�J������P�ы�8�B�PWj�������h�&Q�҃���8�P�B<�M��E�|�Ћ�8�Q�RLj�j�������QP�M��ҡ�8�H�A������R�]��Ѓ������Q������R�Ç��P������h'  P�E�}�ݟ  ������8�Q�B<�M��E�~�Ћ�8�Qj�j�VP�BL�M��Ћ�8�Q�J������P�E�}�ы�8�B�P������Q�]��҃���8�P�B<�M��Ѕ�t�M�Q�� ����8�B�P�M�Q�E�m�҃������;�t	P�o�  ��������;ǉ��������������t	P�J�  �������;ǉ�������������ĸ��t	P�%�  ��������������������������E��� ������E���� ��8�H�A��(���R�E� �Ѓ���ȸ���E�����蕮	 3��M�d�    Y_^[�M�3��E� ��]� ��e �e �e �e �e 	f f f !f )f if �e �e �e �e �e �e �e %f -f 7f Af Kf Uf _f | }| �| \~ \ � ;� � �� c� �� +� �� ������������V��V�+ ���    ^�������������U��V��N��W�}t�F+���;�r�� �F��_^]� �̋Q��u3�3Ʌ�����ËA+���3Ʌ�����������������V��V��H ���    ^�������������U��E�M�@���PQ��� ��]� U��E�U��    QR�� ��]� ��U��E�U��    QR�� ��]� ��U��E��|;A}
�I��]� 3�]� �U��M����w3ɍ�    R�ı  ����]Ã��3����s��EP�M��E    �X� h0�M�Q�E�t$�s� ���������U��EVP���y� �t$��^]� ����U��VW�}��;~tmS3�;�~L9~~�~�N��PWQ����;ÉFtB�V;�~��+ʍI���Q�R��SP�K� ��[�~_^]� �F;�t�SP�B�Љ^�^�^[_^]� �������������̋A�@��Ɂ�   v��|�]UU ;�}���Ã��   ��������������U��SW�}����~b�U��|[V�u��|R;�tN�C�:;�D;�@�K�>;�~�;�}��P��������U�C����Q�R�ЍvQ��P��� ��^_[]� ����������U��VW�}��;~tgS3�;�~F9~~�~�N��PWQ����;ÉFt<�N;�~��+����R��SP�� ��[�~_^]� �F;�t�SP�B�Љ^�^�^[_^]� ����U��S�]��V��~Z�U��|SW�}��|J;�tF�F�;�<;�8�N�;�~�;�}��P���7����U�F��    Q��R��P��� ��_^[]� ��U��VW�}��;~teS3�;�~D9~~�~�N��PWQ����;ÉFt:�N;�~��+���R��SP�� ��[�~_^]� �F;�t�SP�B�Љ^�^�^[_^]� ������U��S�]��V��~Z�U��|SW�}��|J;�tF�F�;�<;�8�N�;�~�;�}��P���7����U�F��    Q��R��P��� ��_^[]� ��U��M����w3�Q��  ����]� ���3����s�EP�M��E    �� h0�M�Q�E�t$��� ��������������U��VW�}��;�tE�G��_�F    ��^]� 9F}P�A����N��t�G�F�W�@���PRQ��� ��_��^]� �����U��V��M��|<�F;�}5+���P�APQ�������F��N�V3��I�ʉ�A�A�A�A�A^]� ��V��~ ��$t%�F��tj P��$�F    �F    �F    ^�����������V��~ �%t%�F��tj P�%�F    �F    �F    ^�����������U��VW�}��;�tB�G��_�F    ��^]� 9F}P�a����N��t�G�F�W���PRQ�� ��_��^]� ��������U��V��M��|-�F;�}&+���P�APQ�������F��N�V3��ʉ�A^]� �VW��3�9>t	V谪  ���>�~�~�~�~_^�������������V��~ �%t%�F��tj P�$%�F    �F    �F    ^�����������U��VW�}��;�t@�G��_�F    ��^]� 9F}P�A����N��t�G�F�W��PRQ�� ��_��^]� ����������U��V��M��|*�F;�}#+���P�APQ���j����F��F�N��    ^]� ����V��~ �,%t%�F��tj P�8%�F    �F    �F    ^�����������U��V��~ ��$t%�F��tj P��$�F    �F    �F    �Et	V�m�  ����^]� ���U��V��~ ��$t%�F��tj P��$�F    �F    �F    �Et	V��  ����^]� ���U��V��~ �%t%�F��tj P�%�F    �F    �F    �Et	V�ͫ  ����^]� ���U��V��~ �%t%�F��tj P�$%�F    �F    �F    �Et	V�}�  ����^]� ���U��V��~ �,%t%�F��tj P�8%�F    �F    �F    �Et	V�-�  ����^]� ���U��E9A}P����]� �����������U���VW�}����}
_3�^��]� S�]���  �F;ǋ��ύ�N�ɉU�u(��8�H��0  h@%h@  �҃�[_3�^��]� ��;��j  )^�F�0  �����j j�и   +�������F�ʙ��߉}���WS�� �ȉU�;�u��E�;�u�;�|�;�r��]�Ù9U�|�;�r��M�F�V��Fы���ɉVh@%u��8�Q���  hV  P�у����8�RhW  PQ��  �у���������V�}���N���F~>+�ɋ�+U��QӍ��Q��P�R� �F+]��    Q��RP�:� ���X  �ɋ�+U�Q��Q��R�� ���9  ��~�V��    Q�R��R��� ���F����V�  �F�D����������؋F���;���   ;���   j jWS�� �ȉU�;��=����E�;��2���;��*���;�� ����E�9U�����;��	������h@%u#��8�Q���  ��    h{  P�у��"��8�Jh|  ��    RP��  �Ѓ����������N���V�^�F9E}"�M�V+���P��P�Eȍ�Q��� ���}�} t=�F;�}�N��+���R��j R�6� ���E�V��    Q��j P�� ���M��N[_�   ^��]� ���U��V��蕟  �Et	V詧  ����^]� ���������������U��S�]V��9^Ws�� �F�}+�;�s����v^�N��r�V��V���Ur�V��V+�P�E��P+�Q�R�� �F+ǃ��~�Fr�N_� ��^[]� �N� _��^[]� ��U��j�h�+d�    P��SVW�  3�P�E�d�    �e����}�E�������v���"�_������������;�s�����+�;�w�4�NQ���E�    �[����E�(�E�M�E���e�P�E��=����E��� Ë}�u�]��v �r�G��GSP�E�VRP�� ���r�OQ�(�  �����M�G�  ��w�_r��� �M�d�    Y_^[��]� �u�~r�VR��  ��j �F   �F    j �F �� �����U���SV��F;FW�}��   �@��Ɂ�   v��|�]UU ;�}�ȍ����   ~� �F����   ��+ȸ���*���������xy;F}t�M�� 9^��G�O�U�W�E�G�M��O�U�E��M�}S�������F�M�@�F�Љ�U�P�M��H�U�P�M��H�U�_�P�F^[��]� 9^}S���k����F�N��@����O�H�W�P�O�H�W�P�O_�H�F^[��]� U��S�]V��FW�~;�ur��    ��   v��|�  ;�}�������   ~� �V��t/��+���x&;�}";��}Q���	����V�F���F_^[]� ;�}Q��������N��V_���F^[]� ���U��E�U+���V�u��    +��~QRQV�� ����^]�U��j�h�+d�    PQV�  3�P�E�d�    h&jhD�j�I�  �����u�3�;��E�t���A�  ��%�ƋM�d�    Y^��]����������V��~r�FP�>�  ��3��F   �F�F^����������̃y$r�AÍA���V��F��t	P� �  ���F    �F    �F    ^�������U��S�]VW�}9_��s��� ��E+�;�s���M;�uj��W������Sj ������_��^[]� ���v�P� �M�F;�s�FPW���t����M��vj�yr/�I�-��u���~r�F_�  ��^[]� �F_�  ��^[]� ���~�^r���ËUW�Q�NQP��� ���~�~r��; _��^[]� ����������U��SV��N��W�^r���ËU;�r1��r���Ë~�;�v��r��EP+�RV�������_^[]� �}���v�X� �U�F;�s�NQW���|����U��vC�N��r����u���~r�_��^� []� ��WRQP�� ���~�~r��; _��^[]� ���������U��E�M�U+�����    V�4tPQPR�N� ����^]� ���������������U��V�u��W�}�Ƌ�v�US��������w�[��_^]� �U��j�h(,d�    PQV�  3�P�E�d�    ��u��+� 3��N��&j��A�A   P�E��A�EP�{����ƋM�d�    Y^��]� �������V����&�~$r�FP�(�  ��3��F$   �F �F��^�n� ��������������U��UV���W�F   �F    �F �x�����u�+�PR�������_��^]� ���U��j�hX,d�    P��D�  3�P�E�d�    jh�&�M��E�   �E�    �E� �����E�P�M��E�    ����h��M�Q�E��&�<� ��U��j�h�,d�    PQVW�  3�P�E�d�    ��u��}W�%� 3�j��N��&�GR�A   �QP�U��Q�����ƋM�d�    Y_^��]� �U��EVP��������&��^]� ����U��j�h�,d�    P��D�  3�P�E�d�    jh�&�M��E�   �E�    �E� �����E�P�M��E�    ����h��M�Q�E��&�<� ��U��j�h�,d�    P��D�  3�P�E�d�    jh�&�M��E�   �E�    �E� �����E�P�M��E�    �G���h��M�Q�E��&��� ��U��SV3�W�};���^�^�^tB�����?v�����SW���������;��N�F�F�ϋ�v�]��������w���V_^[]� �������������U��Q�ESV���M�N��Wu3���~+����]����  ��u3���F+�������?+�;�s�a�����u3���F+����;���   �������?+�;�s3�����u3���F+����;�s��u3���~+����j W������N��P�E�EPQ�������URSP�������MP�FPQ���o����F��u3���N+���م�t	P�p�  ���E����_�V�N�F^[��]� �F�}��+���;Ӎ�    �E��MsG�QPW�������F��+׍MQ��+�SP���/����EF�v�MQ+�VW�M  ��_^[��]� P��+�PS�������U�RSW�F������M�EP�QW�qM  ��_^[��]� �����U��Q�ESV���M�N��Wu3���~+����]����  ��u3���F+�������?+�;�s������u3���F+����;���   �������?+�;�s3�����u3���F+����;�s��u3���~+����j W�"����N��P�E�EPQ��������URSP��������MP�FPQ�������F��u3���N+���م�t	P谚  ���E����_�V�N�F^[��]� �F�}��+���;Ӎ�    �E��MsG�QPW���H����F��+׍MQ��+�SP���o����EF�v�MQ+�VW��K  ��_^[��]� P��+�PS��������U�RSW�F�!����M�EP�QW�K  ��_^[��]� �����U��QSV��W�~��t�F��+���u3��!;�v�� �E��t;�t�� �]+����U�E�MRjPQ���*����~;~v�g� �}�<�;~w;~s�R� �E�x_�0^[��]� �������U��QSV��W�~��t�F��+���u3��!;�v�� �E��t;�t�� �]+����U�E�MRjPQ���Z����~;~v��� �}�<�;~w;~s��� �E�x_�0^[��]� �������U���V��V��u3���N+�����t#�F+���;�s�F�M�����F^��]� W�~;�v�Z� �EPWV�M�Q������_^��]� �������U���V��V��u3���N+�����t#�F+���;�s�F�M�����F^��]� W�~;�v��� �EPWV�M�Q������_^��]� �������U��V�u�F��F������������������� ����������D�Ez��^�P�P�]��������������N�X�N^�X]���U��M�Q���VW�y�I;׍I�Ru3�u�֍֍@�$ƍ��B���`�B�`�� �A�`�A�`�8�4@�E�Ѝ��$��4��B�f�B��f���ȍ��"�@�b�@�b���u�̍U���R��V���]������������]��������]��������_��^��]�����������V����t}��8���   �B4���Ѕ�ui��8���   �B(���Ѕ�uR��8���   �B0���Ћ���t7�I ��8���   �B(���Ѕ�u;�t��8���   �B0���Ћ���u�3�^���������V����t}��8���   �B4���Ѕ�ui��8���   �B(���Ѕ�uR��8���   �B0���Ћ���t7�I ��8���   �B(���Ѕ�u;�t��8���   �B0���Ћ���u�3�^���������U��j�hJ-d�    P�� SVW�  3�P�E�d�    �}3�;ˉ]�u���% �ǋM�d�    Y_^[��]��� ��;��  ��8���   �B����=�  �   �]ԉ]�h�  �M��E�   ��  �   �M��M�S�M�QP���#- ��t&��8���   �PL�M�Q�҃����  ���]�u�E��   �M�u��]��b�  8]�t7���f ��8���   ��U�R�u�]��Ѓ��ǋM�d�    Y_^[��]Ë�8���   �JL�E�P�у�P���� ��8���   ��M�Q�u�]��҃��ǋM�d�    Y_^[��]Ë��� �ǋM�d�    Y_^[��]�����������V����t@���$    ��8�HH���   j h�  V�҃���u��8���   �B0���Ћ���u�3�^�j ���2 ^�����������U���8�H@�U�A,R�Ћ�8�Q��j �ȋB4h�  �и   ]� ���������U��SV�uW��3��9  ��~8�]��$    �N��t�F+���;�r�� �F;�t�΃���8  ;�|�_^3�[]�_^�   []��U��j�hj.d�    P���  SVW�  3�P�E�d�    �ك}�}�5  ��8�H�A�U�R3��Ћ�8�Q�J�E�P�u��эUR�E�P�M�QV�E�舤  ����t#����} u�UR�E�P�M�QV�e�  ����u�j ��腸  ��8�8�  �B��  �P�M�Q�ҡ�8�H�Aj j��U�h&R�Ћ�8�Q�J��d���P�E��ы�8�B�Pj j���d���h&Q�ҍE�P��d���Q��8���R�E��V���M�QP��(���R�E��vV����@P��H����E��� ��h�%�������E��} ��������P�E��k WP�����Q�E��y VP��H���R�E�	�g ��������E��� �������E��� �������E��� ��H����E��� ��8�H�A��(���R�E��Ћ�8�Q�J��8���P�E��ы�8�B�P��d���Q�E��ҡ�8�H�A�U�R�E��Ѓ��1 �Eh1D4ChCD4Cjjj��H���Q��Ȉ]��K ��j hd(��   �M��O��j h�%�M��E��O���U�R��H����E�� P�E�P��t���Q�E���T���U�RP�E�P�E���T��P�E��}�  ��8�Q�J�E�P�E��ы�8�B�P��t���Q�E��ҡ�8�H�A�U�R�E��Ћ�8�Q�J�E�P�E��ы�8�B�P�M�Q�]��҃�0�}  �M��>N��j h�%�M��E��+N��h�%��,����E��g  ��h�%��d����E��Q  ��������P�E��? WP������Q�E��M VP������R�E��; ���M�Q���E�� P�U�R��t���P�E� ��S���M�QP�U�R�E�!�S��P�E�"�H�  ��8�H�A�U�R�E�!�Ћ�8�Q�J��t���P�E� ���E���8�B�P�M�Q�҃�(�������E��B  �������E��3  �������E��$  ��d����E��  ��,����E��  ��8�H�A�U�R�E��Ћ�8�Q�J�E�P�]��у��UR�E�� ����H����E    �E���  ��8�H�A�U�R�E� �Ћ�8�Q�J�E�P�E������у��   �M�d�    Y_^[��]� �P�M�Q�E� �ҡ�8�H�A�U�R�E������Ѓ��M�UWQR��衭  �M�d�    Y_^[��]� �������������U��j�h�.d�    P��0V�  3�P�E�d�    h'  ��u  ���8�H�A�U�R�Ћ�8�Q�J�E�PV�ы�8�B�P�M�Q�E�    �ҡ�8�H�Aj j��U�h�(R�Ћ�8�Q�J�E�P�E��ы�8�B�Pj j��M�h�(Q��j �E�P�M�Qh j �U�RhT� �E���^ ���8�H�A�U��TR�E��Ћ�8�Q�J�E�P�E� �ы�8�E������B�P�M�Q�҃��ƋM�d�    Y^��]������U��j�h�.d�    P��VW�  3�P�E�d�    ����X  �LE  ���E�N�F��M��&� ��8���   �Bx����P�MQ��0  ��P�N �E�    �F� �M�E�����藄 �UR���  ���Et=�EP�M�Q�M�EC  �8 �Eu�B� �E��H;Ju�0� �E�P�B�F(��F(   ���:������K�E���M�t�MQ�U�R����B  �8�@�E���K�M�t;�t��� �U�9U�t)��u��� �E�;Gu�� �M�Q�M�j�V0��� �M�d�    Y_^��]����������������U��j�h./d�    P��   SVW�  3�P�E�d�    �u����  ��8���   �B����=�  ��  �M��(  �C  ��8���   �؋Bx����P�M�Q�p/  ��P�K�E�    轊 �M��E������� ��8�BH�P,������Q�����E�����   �$��4�����4����P�M�Q�/.  ��P���$% ��8�BH�P,������Q�M���E�����   �$��4�����|����P�M�Q��-  ��P���	% 3��}܉}��E�   �}��}�h�_ �M��E���  �uW�U�RP���E��o! �M��E���  h�_ �M�趻  W�M�QP���E��E! �M��E�蹭  ��8���   �P8�M�Q�҃���t_��8���   �A@�U�R��P�MQ��-  ���R����# ��8P���e4 ��8���   �J@�E�P��P�UR�-  � ��P�A��8Q���# ��8���   �P@�M�Q��P�EP�a-  ���Q���4 ��8R���# �}̉}�h�_ �M��E�迺  W�M�QP���E��N  �M��E��¬  ��8���   �P<�M�Q��Q���$�' �}��}�h�_ �M��E��k�  W�M�QP���E��� �M��E��n�  ��8���   �P8�M�Q�҃���wF�$��� j�4��(�����$��! ��(�����$�! j	�
j�j�j���! ���   �� ��8���   �Bx����P�MQ�t,  ��P���   �E�	��� �M�E��� ��   ��8���   ��M�Q�E��ҡ�8���   ��U�R�E��Ћ�8���   �
�E�P�E��ы�8���   ��M�Q�E������҃��   �M�d�    Y_^[��]�3��M�d�    Y_^[��]ÍI �� �� �� �� �� �� �� �� �� ��������U��j�h_/d�    P��|SVW�  3�P�E�d�    ��8�HH�u���   h�  V�ҋ���8�HH��p  3�Sh�  V�}��҉E��8�HH���   h�  V�]��҃��M�QP��x����T  �]�;���|�����   �}�U����U���I �ۋw�t�E�+���;�r�b� ���ۋw�t�E�+���;�r�F� ���ۋ7t�E�+���;�r�+� ���ۋwt�E�+���;�r�� �����m�u��}3��ۉu�u3���E�+���;���  ��t�E�+���;�r��� �<���  ��t�E�+���;�r�� �<�~P�W��u3���O+�����t�G+���;�s�G�0���G� �w;�v�l� �E�PVW�M�Q���AS  �u�3�3�3��M��E��U�3�9]��E��U�]���  �}������}�9>uB�E���t��+�+�����;�s����E���   ;ȋ�v��� �U�R�E�VP�E�P�   9~u5�E���t��+�+�����;�s����E��   ;ȋ�v�� �U��l9~u2�E���t��+�+�����;�s
����E��Z;ȋ�v�u� �U��59~uK�E���t��+�+�����;�s
����E��#;ȋ�v�>� �U��M�QV�E�PR�M��R  �E��M��U���;]��]�������U���%  3ۅ�u3����+���;���  ���E�    t��+���;�r��� �E��M��ɍ<�t��+���;�r�� �E��M��ɍ4�t	+���;�r�� �M�����P�E����T��R��MR�z5 �M�QP�0�������t�E�   �E���t�M���+���;�r�B� �M��E����<�t��+���;�r�%� �M��E����4�t	+���;�r�
� �E���M��R����T
���LRQ�M��4 �U�RP��������t�E��E���t�M���+���;�r赿 �M��E����<�t��+���;�r蘿 �M��E����4�t	+���;�r�}� �E�����Q�M����T
���LRQ�M�]4 �U�RP��������t�E��E���t�M���+���;�r�(� �M��E����<�t��+���;�r�� �M��E����4�t	+���;�r�� �E�����Q�M����
���LRQ�M��3 �U�RP��������t�E��}�t�E��M��������}�W��u3���O+�����t�G+���;�s�G�M�����G��w;�v�`� �U�RVW�E�P���5O  �M��E���u3��+���;���   �}�W��u3���O+�����t�G+���;�s�G�M�����G��   �w;�v�� �U�RVW�E�P�   ��uM�]�S��u3���K+�����t�C+���;�s�C�8���C�m�s;�v蜽 �M�QVS�U�R���N�}�u��W��u3���O+�����t�G+���;�s�G�0���G��w;�v�L� �E�PVW�M�Q���!N  �M�3�;��E� t	Q�N  ���}��|����u��u��u��u���������t	S�$  ���   �M�d�    Y_^[��]�����������U��j�h�/d�    P��|  SVW�  3�P�E�d�    �]3�;���  ��8���   �B����=�  ��  ��8�QH���   h�  S�Ѓ����q  ��8�QH���   VhO  S�Ѓ�;Ɖu��  ���|" ��8�QH�����   h�  S�Ћ�8�Q���  hp(�@��h�   P�ы�8�E�BH���   h�  S�u��у�����   ����    �x&�֋Ǿ   �H��M��H��E��M�������]��E��M��M��������]��E����]��E��]��E�}��]��E��9�}��]؉y�}؉yu��E��؋��8���BH���   h�  S�у�9E��e����
���<9 �E��8�BH���   j h'  S��h�  �E��#{  �����u�3�;��E�tF��8�BH���   h�  S�ы�8���BH���   h�  S�у��}� ����RjWP�\: ���E��E�������  ��8�HH��p  j h�  S�҉E��8�PH�R,����x���P���ҋ��8�   ������j �HH��p  h�  S�ҋM��U��E�}��QR�U���������$QRPW��8����S  ��8�HH���   h�  S�E�   3��҃�����   �}���3�;G�U���Rj V�E�    �M؍�8����*K  �E�PjV��8����K  �M�QjV��8����K  �}� ��   �U�RjV��8�����J  �U�E��M܉U��U��EĉMȉŰM�E�P���+  ��8�QH���   h�  S�����Ѓ�;��K����}�}� t�M�Q��w  ����Bj ���Ѕ�t~�M�U�]WQ�MR�U�������<������P��8���QR��V�E�P�E������C  ��<���Q��z  ���   �M�d�    Y_^[��]ËE��M܉E��E��MĉẺE��'�����Bj���Ћ�8�Q�J�E�P�ы�8�B�Pj j��M�hH)Q�ҍE�P�E�褃  ��8�Q�J�E�P�E��ы�<������P��8���QR��V�U�R�E�������B  ��<���P�z  ��3��M�d�    Y_^[��]�����U���8�HH���   S�]VWS�ҋu(�}����t)�M$�E�UVQ�M���$R�UQWPR������$��   ��8�HH���   j S�ҋM�؃���tH��8���   �B��=__ t=�  t�M$VQ�VP�E�U�E�M���$RPWSQ�N�����$�p��8�B@�PQ�҃��   uW��8���   �]�B����-�  t��u6�E���$��WQ�M�������E�U�E�M���$RPWSQ���������8���   �M�P4�ҋ؅���   ��tR��8���   �M�B��=__ t	�}$__ u/��8���   �M�BV���E�M�UP�E���$QRWSP��M$�E�U�EVQ�M���$RPWSQ�D�����$��t3���8���   �P(���ҋ؅��c���_^[]����������U��j�h�1d�    P��	  �  3ŉE�SVWP�E�d�    �M�E�}�����3���������x����������������$� �������u����	 h'  �,`  P������R��  ��P��t����E��x �������E� �mp h'  ��_  P������P�  ��P��x����E���w �������E� �4p h'  �_  P������Q�]  ��P��|����E��w �������E� ��o ��8�B@�H,W�у�h��hE  ����E �����R��,���Q���
 ����������	wM�$��� �   �A�   �:�   �3�   �,�   �%�   ��
   ��   ��	   �	�   �3�P��(������ ݅,�����ݝd����G�  ��;���  ���$    �d$ ��8���   �P����=�  �j  ��H����G.  ���ω������� ���Q$ +�t	��uj�j���� ��8���   �Bx����P������Q��  ��������P��X  �E��Cv �������E� �n ��8�BH�P,������Q����݅d������$����4����   �������݅����P���������\$݅ ����\$݅�����$�0� ���	� ��4���Q�������g� ��8�BH�P,������Q����݅d������$����4����   ��P����݅����P���������\$݅�����\$݅�����$�� ���� ��������4���Q��訤 h(����<� ���  ���O� �    �hY����" ��ݝ�����o# ��$��������ܽ�����*�$茑 3���T�����\���h�  ��L����E�誦  V��T���RP���E��6 ��L����E�觘  ��8���   �A<��T���R��ݝ������8�QH�R,��������P���ҹ   ���������݅����������܅����݅��������݅����݅��������݅������܅����݅����������܍������݅�������̍�4���������܅����݅����������܍������݅d����$P���\$���\$�$�� ����� ��4�����8������ĉ��<����P��@����H��D����P��H����H�������P�� ��8���   ���T���R�E� �Ѓ�3�3����������;��e�����������!  �������@�������@������� �������@�������������E��q�  ��;���  ��$    ��������(  �؋��LY ��8���   �Bx����P������Q�L  ��P�K�E��r �������E���j ������������P��`���Q�������������������b?  ��8���   �P����=G  ��  ��T�����\�����8�HT�QVW�E�	�҃���t6h4  ��L������  ������V��T���QP���E�
�	 ��ƅ����uƅ���� �������E�	   t���������L����ϕ  ������ �c  ��8���   �P@��T���Q�҃����������S �F���\$�������F�\$��$�iV �������C(�C$��8�HT�Qj W�ҍ�l���Q�����������l����E����  ����   ������:�  ��������������R�E��R�  ��l���QV��RP�E��{  �����������E����  ������E����  ��tf��<���P��l�����  P������Q�E��C  ��j���E��Ck P���\ �������E���h ��8�B�P��<���Q�E��҃���l����E�	�a�  ���8�C(��8�K$��8�BT�HjW�у���t7h�  ��4�����  ������j ��T���RP���E�� ��ƅ����uƅ���� �������E�	   t���������4����֓  ������ tS��8���   �A@��T���R�Ѓ����������Q �F���\$�������F�\$��$�uT �������K,�	��8�S,��8�HT�QjW�҃���u��8���[P�C0��8�QT�BjW�Ѓ�����  3��u��u艵����������$�����,���h`	  ��D����E��ݠ  V�M�QP���E��l ��D����E��ݒ  ha	  �����譠  V�����RP���E��9 ������E�誒  h�  ��l����z�  V��$���QP���E�� ��l����E��w�  ��8���   �P@�M�Q�҃����������RP �F���\$�������F�\$��$�!S �������C8��8���   �J<�����P���[X��8���   �P<��$���Q���[@��8���   ���$���R�E��Ћ�8���   �
�����P�E��ы�8���   ��M�Q�E�	�҃�����[X��8�HT�QjW�ҡ�8�HT�QjW�ҡ�8���   ���T���R�E��Ѓ�3���8���   �B(���Ћ�;��O�����������  ����������������  �������@�������@������� �������@������;��E���  ��8���   �BX���Ѕ��v  ������������R��`���������P��������������8  ��8���   �BX���Ћ�;��  ���    ������������R��`���������P�������������8  �������"  ����葄 ��8���   �Bx����P������Q�  ��P�Oh�E��l �������E��Rd ������j R���  ���~ ����P��� �~ ��Q���� ��������M �F8���\$�������F0�\$�F(�$�P ������R���g� ��W�.~ ��3��������؅��������8���   �������BX�Ћ����������d  ����8���   �B0���Ѕ���������   ������Q��l���R�������6"  ���> u�4� ��N;Hu�%� �V�B������k�p�T�|�\�D�@�������U�Q�����R�������E���!  ���> u�ا ��N;Hu�ɧ �V�B������k�p�U苵�����D�M�8�X�P�H3����������������������l�������   h'  ���#R  P������R��  ��P�Oh�E��j �������E��gb j���� V���6� VVV�������O � P��较 ���������1�  ����te�	��$    ����8���   �Bj����݅d���P���$������Q������R������PVW�������8���   �B(��$���Ћ���u���8�Q@��x����J,P�ы�8�R��j �ȋ��   h�  �Ѕ���  ��腺  �؅ۉ�������  ��I ��8���   �B����=�  �m  ��8�QH�R,������P���ҋ�   ���������e ��3�����  ��8�HH��p  Wh�  S�҉�x�����8�HH��p  Wh(  S�ҋ��8�HH���   h(  S�������������҃� ����  �ލI hp(h  hD�j,�Zh  �����������E�t�Qjj j����< ���3��; �E�ǅ����    ~y�������@��x����|�݅d������$�������G�Q���\$��p�����\$�G��$�� ����� ������������RP��� ����������;������|�����$��j �� 3�9������~-���$    �ۅ�������x���$W� ��;������|݋������ۅ���������$P���~ ��Bj ���Ѕ�tX�������  ���w���8���   �������Bx��P��P���Q�x  ��P�O �E���f ��P����E��_ �]��8�B�P�M�Q�ҡ�8�H�Aj j��U�h *R�ЍM�Q�E��o  ��8�B�P�M�Q�E��ҋ�P��j���ҋ��8������������QH���������   h(  ��P���������у�;�������������  ;��N  ��8�BH��p  Wh�  S�ы�8W�������BH��p  h(  S�ы�8���BH���   h(  S�������������у� ���  �����$    �d$ hp(ho  hD�j,�e  ����x������E�t����	 ���3��G(   �; �E�ǅ����    �   �������@�������t��	��$    ���F���܍����������܅�����F�܍������݅��������F�܍����܅�����F�܍������݅��������F�܍����܅�����F�܍������݅�������݅d����$Q�����\$��p����\$�$��� ���� ������R�O����ۅ�����{ t�3������x���ۅx�������t���ݝt���Q�O�  ����������;������������{ ��   ������݅�����@�������ЍЃ�������܅�����@܍������݅�����H��݅�����܅�����@܍������݅�����H��݅�����܅�����@܍������݅�����H��݅d����$Q�����\$��p����\$�$��� ���� ������R�O�����荅l���ݝl���P�O�  ��Bj ���Ѕ���   �������  ���N�~�輸 ��8���   �������Bx����P������Q�  ��P�N �E���b �������E��'[ ������R���)�  ����x�����   ��x���P�����Q��������  ���? u��� ��G;Bu豟 �O�Q�V(�h��8�H�A�����R�Ћ�8�Q�Jj j������h�)P�э����R�E���j  ��8�H�A�����R�E��Ћ�B��j���Ћ��8������������BH���������   h(  ��Q���������҃�;��2����������2  ��8�H�A��T���R�Ћ�8�Q�JWj���T���h�)P�ы�8�B�P��$���Q�E� �ҡ�8�H�AWj���$���h�)R�Ѝ�<���VQ�E�!�01��P��$���R��\���P�E�"�H%����T���QP��<���R�E�#�0%����HP�E�$�i  ��8�H�A��<���R�E�#�Ћ�8�Q�J��\���P�E�"�ы�8�B�P��<���Q�E�!���E� ��8�H�A��$���R�Ћ�8�Q�J��T���P�E��у�3��������؅ۉ������\���j<��i  ���������'� jA��i  ����|����Y hp(h�  hD�j<�L`  ��������3�;��E�&t��|���R���h	 �������������9������E�%��   ��|����E��>X �������P������QR��W��l���P�E��(  ������Q�_  ��������P������Q�������������R��W��l���R�E� �;)  ������P��^  ���������������������E�����螺 ������  ��L���Q�������  ��8�B�PdV��L����E�'��hp(��h�  �ChD�P�`  ����8�P��V�CP�BhW��L����Ћ�����QVjW������� �G{ �؄�uQ��8�B�P�M�Q�ҡ�8�H�AVj��U�h�)R�ЍM�Q�E�(�)g  ��8�B�P�M�Q�E�'�҃�;�t	W�^  ��jd��g  ��|���P��<���Q�1��P�E�)��f  ��8�B�P��<���Q�E�'�ҋ���������j�҄��E�%��   ��8�H�A��L���R�Ѓ���|����E��CV �������P������Q��RW��l���Q���E��&  ������R�]  ��������P������Q�������������R��W��l���P�]��?'  ������Q��\  ���������������������E�����袸 ������   ��8�B�P��L���Q�҃���|����E��U �������P������QR��W��l���P�E���%  ������Q�Q\  ��������P������Q�������������R��W��l���R�E� �~&  ������P�\  ���������������������E������� 3��M�d�    Y_^[�M�3��q� ��]� ��� �� �� �� �� �� �� �� �� �� ��������U���E�E��V�u���$V�@���\$�M��@�\$� �$�k� ���D� ��^��]��������������U���E�E��V�u���$V�@���\$�M��@�\$� �$�� ����� ��^��]��������������U��V�u���= �E�@���\$���@�\$� �$�r@ ��^]��������������U��Q��8�P�M�BdSVWj �E�    ��h�'��h  �_hD�S�6\  ��8�Q�M��j ���BhSV���> �}V���Z ��t	V�Z  ����_^[��]�������̋Q��u3�ËA+�����������������U��E��y u������y t�]�����U��U�BV�0�r�0�~ u�V�r�p�I;Q^u�A��B]� �J;u���B]� �A��B]� �������������U��U�V�p�2�p�~ u�V�r�p�I;Q^u�A�P�B]� �J;Qu�A�P�B]� ��P�B]� ���������U��E�H�y u����H�y t�]����U��E�H�y u����H�y t�]����U��E��y u������y t�]�����V��> u譖 �F�x t^鞖 �H�y u��x u�I �ȋ�x t��N^Ë@�x u�N;Hu�F�ЋB�x t�F^��������������U��VW�}��;~tfS3�;�~E9~~�~�N��PWQ����;ÉFt;�N;�~��+���R���SQ�b� ��[�~_^]� �F;�t�SP�B�Љ^�^�^[_^]� ����̋A��    ��   v��|�  ;�}���Ã��   ����������������U��j�h!2d�    PQ�  3�P�E�d�    �M�M����E�    t��� �M�d�    Y��]� ������U��j�hQ2d�    PQ�  3�P�E�d�    �M�M����E�    t�w? �M�d�    Y��]� ������U��j�h�2d�    PQ�  3�P�E�d�    �M�M����E�    t��� �M�d�    Y��]� ������U��j�h�2d�    PQ�  3�P�E�d�    �M�M����E�    t�'& �M�d�    Y��]� ������U��j�h�2d�    PQ�  3�P�E�d�    �M�M����E�    t�g( �M�d�    Y��]� ������V��> u�� �F�x t^�ޓ �H�y u��x u�I �ȋ�x t��N^Ë@�x u�N;Hu�F�ЋB�x t�F^��������������U��U�BV�0�r�0�~ u�V�r�p�I;Q^u�A��B]� �J;u���B]� �A��B]� �������������U��U�V�p�2�p�~ u�V�r�p�I;Q^u�A�P�B]� �J;Qu�A�P�B]� ��P�B]� ���������V��> u轒 �F�x t�@�F�x te^颒 ��y u �A�x u��$    �ȋA�x t��N^Ë@�x u��$    �N;u�F�ЋB�x t�N�y t^�F� �F^��������U��E9A}P�?���]� �����������U��S�]��VW��}W�~ tB�~��x$��iۘ   �N��P�j �҃���   ��}�N��Pj Q�����F    3�_�F�F^[]� �F;��~   �N��PSQ����3�;FtZ�N��+�iɘ   i��   WR�Q�ڑ �F��;�})����i��   +ȉM��F�P�������ǘ   �mu�_�^^[]� _�V�V^[]� ~a���;�|2��+�i��   ���E��$    �N�9�B�j �Ё�   �mu�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^[]� ������U��S�]��VW��}Q�~ t<�~��x��k�p�N��P�j �҃���p��}�N��Pj Q�����F    3�_�F�F^[]� �F;�}u�N��PSQ����3�;FtQ�N��+�k�pk�pWR�Q芐 �F��;�}&����k�p+ȉM�d$ �F�P��������p�mu�_�^^[]� _�V�V^[]� ~T���;�|%��+�k�p���E�N�9�B�j �Ѓ�p�mu�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^[]� ������V��> u�m� ��N;Hu�^� �F��^�������������U��j�fO  ����t)�M�U��M�H�M�P��P�I�U�H�P�@ ]� ��j�)O  ����t�     �H��t�    �H��t�    �@�@ ����������U��j��N  ����t/�M�U��M�H�M�P��P�Q�P�I�U�H�P�@ ]� ������������j�N  ����t�     �H��t�    �H��t�    �@�@ ����������U��SVW�}� �ً�u�FP��������6W�:P  ���~ ��t�_^[]� ��������U��SVW�}� �ً�u�FP��������6W��O  ���~ ��t�_^[]� ��������U���SV��F�V;�W�}��   ������   v��|� � ;�}�������   ���^��tQ��+���xH;�}D;ЋO��M�O��M�}P��������F�U�M���F��P�H�x�F_^[��]� ;�}P��������F���F��O�H�W�P�O_�H�F^[��]� �����U���S�]V��FW�~;�uz��    ��   v��|�  ;�}�������   ~� �V��t7��+���x.;�}*;���]�}Q��胜���V�E��F_�ЃF^[��]� ;�}Q���^����N��V_�ʃF^[��]� ������U��E�M;�t�UV�2�0��;�u�^]��U��SVW�}����}R�~ t=�~��x��i�(  �N��� ����(  ��}�N��Pj Q�����F    3�_�F�F^[]� �F;�}}�N��PWQ����3�;FtY�N��+�i�(  i�(  SR�Q�Ӌ �F��;�}(�؋�i�(  +ȉM�F�P��������(  �mu�~_^[]� _�V�V^[]� ~V���;�|'��+�i�(  ���E��N��� ��(  �mu�9~~�~��F�RWP�Ή~��3�;��Fu�N�N_^[]� �����������U��SVW�}����}R�~ t=�~��x��iې  �N�� ����  ��}�N��Pj Q�����F    3�_�F�F^[]� �F;�}}�N��PWQ����3�;FtY�N��+�iɐ  iې  SR�Q胊 �F��;�}(�؋�iې  +ȉM�F�P���]����Ð  �mu�~_^[]� _�V�V^[]� ~V���;�|'��+�iې  ���E��N��� ��  �mu�9~~�~��F�RWP�Ή~��3�;��Fu�N�N_^[]� �����������U��SVW�}����}P�~ t;�~��x����N��" �����   ��}�N��Pj Q�����F    3�_�F�F^[]� �F;�}{�N��PWQ����3�;ÉFtW�V��+ʍI�R��Q���SR�5� �F��;�}&�@����+ȉM�F�P���a������   �mu�~_^[]� _�^�^^[]� ~Z���;�|+�@+������E��$    �N��F ���   �mu�9~~�~��F�RWP�Ή~��3�;��Fu�N�N_^[]� �����������U��j�h3d�    PQV�  3�P�E�d�    hp(jhD�j��J  �����u�3�;��E�t����A  �(�ƋM�d�    Y^��]����������U��Q�B�x VW�}u�7;p}�Ћ ��@�x t�q�F�x u�?9x}�@���� �x t�E_�p��H�P^]� V��F�V;�u@��iɘ   ��   v��|�Ky ;�}�������   ��;�}2P��������(i��   Fj ��ȋB�ЋNiɘ   NQ�������N��i��   F���N^������V��F�V;�uN��k�p��   v��|�,I ;�}�������   ��;�}=P�������N��k�pF���N^�k�pFj ��ȋB�ЋNk�pNQ���S����N��k�pF���N^�U��E9A}P����]� �����������U��Q�B���x VW�}u�7��$    9ps�@��Ћ �x t�A;ЉU��M�t�7;rr�M��	�M��E�M���E�I_��H^��]� �����V��N�V;�u>��i�(  =   v��|��� ;�}�������   ~�	;�},P���G����"i�(  N��� �Ni�(  NQ�������N��i�(  F���N^��������������V��N�V;�u>��i��  =   v��|�� ;�}�������   ~�	;�},P�������"iɐ  N�� �Niɐ  NQ�������N��i��  F���N^��������������V��F�V�@��;�uJ��   v��|���
 ;�}�������   ��;�}8P��������N�I��F���N^�N�� �F�@��V��R�����N�I��F���N^����U��V����&�~$r�FP��E  ��3��F$   �F �ΈF�<� �Et	V��E  ����^]� ������U��j�hH3d�    P��DSVW�  3�P�E�d�    ���TUUrCj3�h�(�M��E�   �u��E� �~����E�P�M��u�诤��h��M�Q�E��&�4� �U�G�uj RPVP�F����ȋG�   _;��Mu�H�G��W�J�!�} t��G;0u���N�G;pu�H�Q�z �A����   ��Q;
uN�R�z u�Y�Z��J�A ��r�y;qu
��V�������F�X�N�Q�B �F�HQ��������J��z u�Y�Z��J�A ��r�,;1u
��V�������F�X�N�Q�B �F�HQ���>����V�z �F�O����M�G�P�E�Z�H�8�M�d�    Y_^[��]� ������U��j�hx3d�    P��D�  3�P�E�d�    jh�&�M��E�   �E�    �E� �ʡ���E�P�M��E�    �����h��M�Q�E��&�|� ��U��j�h�3d�    P��PSVW�  3�P�E�d�    �M��E�x tCj3�h )�M��E�   �u��E� �M����E�P�M��u��~���h8%�M�Q�E��(�� �؍M�]��������x t�{��S�z t���
�M;ˋyur� �su�w�M��A9Xu�x�9u�>��~�A9u� t���W�����M����Q��I9Y�M�ux� t�ƉA�kW�A����M���A�Z�H��;Ku���� �qu�w�>�S�Q�C�H�U��B9Xu�H��C9u���H�C�A�S�A�Q�C�E�8X��   �M��Q;z��   8_��   �;�ue�F�x u�XV�F ������F�M��x ut�8Zu�P8Zta�P8Zu��ZP�@ �����F�M��V�P�^�@V�X�����t�x u�XV�F �������M��x u�P8Zu�8Zu�@ �A��;x�v�J����0�8Zu�P�ZP�@ �0�����M��V�P�^� V�X�w����_�M�Q�A  �M��A����v����A�E�U�M��H�M�d�    Y_^[��]� ������U��EVP���q�����(��^]� ����U��j�h�3d�    P��PSVW�  3�P�E�d�    �M��E�x tCj3�h )�M��E�   �u��E� �m����E�P�M��u�螟��h8%�M�Q�E��(�#~ �؍M�]��L�����x t�{��S�z t���
�M;ˋyur� �su�w�M��A9Xu�x�9u�>��~�A9u� t���W������M����Q��I9Y�M�ux� t�ƉA�kW�����M���A�Z�H��;Ku���� �qu�w�>�S�Q�C�H�U��B9Xu�H��C9u���H�C�A�S�A�Q�C�E�8X��   �M��Q;z��   8_��   �;�ue�F�x u�XV�F �J����F�M��x ut�8Zu�P8Zta�P8Zu��ZP�@ �x����F�M��V�P�^�@V�X������t�x u�XV�F �H�����M��x u�P8Zu�8Zu�@ �A��;x�v�J����0�8Zu�P�ZP�@ ������M��V�P�^� V�X������_�M�Q�+>  �M��A����v����A�E�U�M��H�M�d�    Y_^[��]� ������U��j�h4d�    P��PSVW�  3�P�E�d�    �M��E�x tCj3�h )�M��E�   �u��E� 譛���E�P�M��u��ޜ��h8%�M�Q�E��(�c{ �؍M�]�������x t�{��S�z t���
�M;ˋyur� �su�w�M��A9Xu�x�9u�>��~�A9u� t���W�
����M����Q��I9Y�M�ux� t�ƉA�kW������M���A�Z�H��;Ku���� �qu�w�>�S�Q�C�H�U��B9Xu�H��C9u���H�C�A�S�A�Q�C�E�8X��   �M��Q;z��   8_��   �;�ue�F�x u�XV�F �����F�M��x ut�8Zu�P8Zta�P8Zu��ZP�@ �����F�M��V�P�^�@V�X�=����t�x u�XV�F ������M��x u�P8Zu�8Zu�@ �A��;x�v�J����0�8Zu�P�ZP�@ �������M��V�P�^� V�X�'����_�M�Q�k;  �M��A����v����A�E�U�M��H�M�d�    Y_^[��]� ������U����Q�B�x S�]V���E�u W�;;x���҈U�t� ��@�x t�_�E�SVP�U�R�$����ȋ�E�I^��H�@[��]� ���������U��j�h84d�    P��DSVW�  3�P�E�d�    ������rCj3�h�(�M��E�   �u��E� �~����E�P�M��u�诙��h��M�Q�E��&�4x �U�G�uj RPVP������ȋG�   _;��Mu�H�G��W�J�!�} t��G;0u���N�G;pu�H�Q�z �A����   ��Q;
uN�R�z u�Y�Z��J�A ��r�y;qu
��V��������F�X�N�Q�B �F�HQ���:����J��z u�Y�Z��J�A ��r�,;1u
��V�������F�X�N�Q�B �F�HQ�������V�z �F�O����M�G�P�E�Z�H�8�M�d�    Y_^[��]� ������U��j�hh4d�    P��DSVW�  3�P�E�d�    ������rCj3�h�(�M��E�   �u��E� 辖���E�P�M��u�����h��M�Q�E��&�tv �U�G�uj RPVP�����ȋG�   _;��Mu�H�G��W�J�!�} t��G;0u���N�G;pu�H�Q�z �A����   ��Q;
uN�R�z u�Y�Z��J�A ��r�y;qu
��V���8����F�X�N�Q�B �F�HQ���z����J��z u�Y�Z��J�A ��r�,;1u
��V���L����F�X�N�Q�B �F�HQ��������V�z �F�O����M�G�P�E�Z�H�8�M�d�    Y_^[��]� ������U���SV��F�W�}���M�t;�t��t �];]�uZ�E���V�U�t;�t��t �E;E�u<�N�QR�������F�@�F�F    � �F�@�F��E_�0^�H[��]� ��t;}t�t ;]t�M����SW�U�R�������]�}�ЋE�8_^�X[��]� ����������U���SV��F�W�}���M�t;�t�'t �];]�uZ�E���V�U�t;�t�	t �E;E�u<�N�QR��������F�@�F�F    � �F�@�F��E_�0^�H[��]� ��t;}t�s ;]t�M�����SW�U�R�������]�}�ЋE�8_^�X[��]� ����������U���SV��F�W�}���M�t;�t�Ws �];]�uZ�E���V�U�t;�t�9s �E;E�u<�N�QR���)����F�@�F�F    � �F�@�F��E_�0^�H[��]� ��t;}t��r ;]t�M� ���SW�U�R�������]�}�ЋE�8_^�X[��]� ����������U��Q�ESV���M�N��Wu3���~+����]����  ��u3���F+�������?+�;�s������u3���F+����;���   �������?+�;�s3�����u3���F+����;�s��u3���~+����j W�B����N��P�E�EPQ�������URSP�������MP�FPQ���ϒ���F��u3���N+���م�t	P��3  ���E����_�V�N�F^[��]� �F�}��+���;Ӎ�    �E��MsG�QPW���h����F��+׍MQ��+�SP��菒���EF�v�MQ+�VW�	�����_^[��]� P��+�PS�������U�RSW�F�A����M�EP�QW�������_^[��]� �����U���S�]VW���w�F�x ��M�u�;P�����ɈM�t� ��@�x t�ɋ։U��}�t:�G;0�M�u(SVjQ��������ȋ�E�I_^��H�@[��]� �����U��B;s�M�SVQ�U�R�E�M�_^��P�@ [��]� ��U���S�]VW���w�F�x ��M�u�;P�����ɈM�t� ��@�x t�ɋ։U��}�t:�G;0�M�u(SVjQ�������ȋ�E�I_^��H�@[��]� ������U��B;s�M�SVQ�U�R�E�M�_^��P�@ [��]� ��U��SV3�W�};���^�^�^tB�����?v����SW�}������;��N�F�F�ϋ�v�]��������w���V_^[]� �������������U��QSV��W�~��t�F��+���u3��!;�v��n �E��t;�t��n �]+����U�E�MRjPQ�������~;~v�n �}�<�;~w;~s�n �E�x_�0^[��]� �������U��j�h�4d�    P���   SVW�  3�P�E�d�    ��E���O  �$��(�E�N����+�E�N���T��E�N���T��E�N���T�E��E�P�M�Q�ΉU��R����8���H�P�X��D�����H���t;�t��m ;�H����k  �}�]��t;�D���t�m ;�H����+  ��u�m ;_u�m �E9C�.  �~ �  ;_u�vm ;_u�lm �K�V���;Cu3��   ;_u�Jm ;_u�@m �K�V���D;Cu�   �V�M������H�V���|�M������;u�   �,�M��{����P�F���M�|�f����;��  �   �U�;Zu��l �C�N���@����U��E��P�@�E��E�U��U���@����P�@�M��e��EĉU��]��E����]��E���'����������  �E��e��]��E����]��E�������A��  �E��e��]��E����]��E�������A��  �~ �~  ��L��������N��  �M�E��w�����8�QD�@��L���Q�J,P�E�P�����U؃����U��]�wa�$��(݅L����]�݅T����]�݅\����=݅d����]�݅l����]�݅t����#݅|����]��E��]��E���E��]��E��]��E��]؋�8�BD�U��L���Q�M�R�P,Q����E�������$��(������݅L���݅T���݅\����=������݅d���݅l���݅t����#������݅|����E��E���������E��E��E����E���������'���������D  �E�������������A�0  �m���������A�"  �M������@�M�}���t;�D���t�mj ;�H�����  �N�Q�E��F8�E�V�@�ʍʃ���4����F �FP�H���Fh�H���F@��F(�FX�H���Fp�H���FH��F0�F`�H���Fx�H�E���݆�   �$P�����\$�\$�$��� ���՚ �}��M�Q�NR�S� ����   �N����   �]��E�����@�$��P�M�Q�_�����N��PR�� ��   �����؍M��m����]�}�����;_u�Ri �K�U�
�����j h)��<����������<���R�E�    �4  ��8�H�A��<���R�E������Ѓ�2��M�d�    Y_^[��]� �FE��NPQ�U�R�n�������$�E�P��4���Q�F�����N��PR�'� �]�N����   ��ݕ\���ݕT���ݕL���ݕt���ݕl���ݕd����U��U�ݕ|����U��U��]��i�  ��8�QD�R,��L���QSP�ҋE����t7��t$��t݅L���݅T���݅\����+�E��E��E�� ݅|����E��E��݅d���݅l���݅t�����]؋N���\$�$P�� �M�?�U�R�E��M�P�Ή}��]�������M�d�    Y_^[��]� �I �!�!""�$�$�$�$
%$%>%R%U���V��F�PVQV�E�P��������NQ�z)  ��3��F�F^��]�����������U���V��F�PVQV�E�P��������NQ�:)  ��3��F�F^��]�����������U��SVW��������E�M�U�u�C�@�C�@�C� �C�@�E�K�M$�C�E �K�C�{ �C    �S�   �ݛ�   _^��[]�  �������U���V��F�PVQV�E�P���S����NQ�(  ��3��F�F^��]�����������U��j�h�4d�    P��VW�  3�P�E�d�    �E�    ��8�P�E�RPP�EP�E�P�ҋ���8�H�u�QV�E�   �ҡ�8�H�QVW�ҡ�8�H�A�U�R�E�   �E� �Ѓ��ƋM�d�    Y_^��]� ������������h'  �F  ����̡�8��t	P�'  ����8    ����U��j�h�5d�    P��  �  3ŉE�SVWP�E�d�    �}�]3��񉅘����������F�$0  ��u�F   3��  ��8�P�B<���Ѕ��v  ��8�Q�Bdj ���Ћ�8�Q�Rhj ��j@��p���P���ҍ������`  ���V��u���P�������E�    �C  ��`���Q�������q  ��u��������  3���5`���R��5p���h0*P��o ������|ۋ�8�E� �Q�J������P�ы�8�B�@j ���V��p���Q������R�Ѓ���8�Q�R|������P���E��҅���8�H�A������R�������E� �Ѓ������� �u�t�������A   �������
  3��2  ��������  ��8�B�Pdj ���ҋ��8�P�Rhj j@�E�P���ҍ�����  ���V�E��   P������}���
  ��L���Q������%
  ����  3��	��$    ����5L���R�D5�h0*P�n ������|ދ�8�E� �Q�J������P�ы�8�B�@j j��M�Q������R�Ѓ���8�Q�R|������P���E��҅���8�H�A������R�������E��Ѓ������� t&�������A   ������E������  3���  ��8�B�P<���҃� ��   ��8�H�A������R�Ћ�8�Q�Jj j�������h(*P�у�jj ��t���R���E�ǅ����   ������8�Q�Rx������Q���E�   ǅ����   �҅�u ��8�H�Q4jS�҃�f=- ƅ����tƅ���� �������   �u�t��8�H�A���������t���R�Ѓ��������}�t��8�Q�J������P�у������� ��   ��8�B�P������Q�ҡ�8�H�Ij j��U�R������P�у�jj��t���R���E�������8�Q�R|������Q���E��҅���8�H�A��t���R���E��Ћ�8�Q�J������P�E��у���t�������r����������E�������   ����M�d�    Y_^[�M�3��#\ ��]� ���U��j�h�5d�    PQV�  3�P�E�d�    h8*h�   hD�j�#  �����u����E�    t���a �*���3Ʌ��E�������8t%jh� �a ��t�   �M�d�    Y^��]�3��M�d�    Y^��]�����������*����������3��A�A�A`�A#Eg�A�����A�ܺ��AvT2�A���ÈAd�Ae�����������̋�3�� �*�H�H�H`�@#Eg�@�����@�ܺ��@vT2�@���ÈHd�He����U���P  SVW�M�3��A!3Ҋp��x�����P�����x���׉������3Ҋp��x��P�����x�����x��������3Ҋp��P�����x�����x��������3Ҋp��P�����x���׃���������m����������E�   �P�3P�X�3X33X�p�x�3�3����ÉX$�X3X��P 3X��3ދp�3p���3�3��ƃm��X�pu��Y�A�Q�q�I�]��M��E�    �I ����#�����#�ϋ}���������M��y�Z�]����u�M�����U���#��#��U�������������y�Z�U����U�U��M�������#Ɖ]�#�Ë]���������E��y�Z�u�u�������#ˉU�#�ʋU�E�����������]��y�Z�U��E����ډu��M���#�#���ދu���������E�E���1�y�Z�u��������ى]��}�������   ����3�3���������]��������n�]��u�M�����3�3���������u�1���n����3ÉU�U�3M�����������E��������n�΋u��]��U��E�����3U���3���������U��������n�E��u��M���3u���3���������u������n�E�E�����(�M��%����E�(   ��M�u���#���#���]�����������ܼ��}��M���M���#��#��]�����������ܼ����U�U��#��E��M���M��#���������E���ܼ����E�E��}����#��M���M��#������������ܼ��u��u��U����#��u��M���#���������u���M�u�ܼ����E����M�����<�]�������<   �}���M��3�3��������}�����bʋ]����M����u�M��3�3�������������bʋ�3ÉU�U��M���M�3�������������bʋ�3ʉu�u�3��������E���E�]���bʋ]����U��U��M���3���M�3�������������bʉE�E�����P�u��M��}��%����}��_ًOȋGU�G�GƉG�G_�O�G�G`    _^[��]������SV��F`W�D0 ��   ~`��7�F`~D�@   2�;�}���    �\0 ~`�F`;�|���{����8   9N`}/��F`�\ ~`9N`|���8   ;�}2ۍd$ �\0 ~`�F`;�|��N�V�F�NX�N�VY�V�N[�N�FZ�F�V\�V�N^_�F]�V_��^[� ���U��V��~e t2�^]� �~d u	�"����Fd�N�E��V�P�N�H�V�P�N�H�^]� �������U��} V��tR�~d uQ�~e uKSW�}�   )]�~e u1�F`��L0 ^`�F�F`u^u�^e��@u���\�����} u�_[^]� �Fe^]� ����U��]�����������U��j�EP�r���]� ��������������U��j�EP�R���]� ��������������U��V�u���W��t�Ej�EP��� ����F����u��_^]� ��������������U��V�u���W��t�Ej�EP��������F����u��_^]� ��������������U��Vj�EP��������^]� ��������U��Vj�EP��������^]� ��������U���EV����*t	V�X  ����^]� ��������������U���8�P�E���   ��VWP�EP�E�P�ҋu����8�H�QV�ҡ�8�H�QVW�ҡ�8�H�A�U�R�Ѓ�_��^��]� ������������U��E��u��8�MP�EPQ�=  ��]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3h�*j;hD�j�-  ����t
W���Ή  �3����Fu_^]� �~ t3�9_��^]� ��8�H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   ��8�H<�Q��3Ʌ����^��������������̃y t�   ËA��uË�8�R<P��JP�у��������U����u��8�H�]� ��8�J<�URP�A�Ѓ�]� ���������������U�졸8��u��8�H�]Ë�8�J<�URP�A�Ѓ�]�U�졸8��$��Vu��8�H�1���8�J<�URP�A�Ѓ�����8�Q�J�E�SP�ы�8�B�P�M�QV�ҡ�8�H�A�U�R�Ћ�8�Q�Jj j��E�h�*P�ы�8�B�@@�� j �M�Q�U�R�M��Ћ�8�Q�J���E�P���у���[t.��8�B�u�HV�ы�8�B�P�M�Q�҃���^��]á�8�P�E��RHjP�M��ҡ�8�P�E�M��RLj�j�PQ�M��ҡ�8�H�u�QV�ҡ�8�H�A�U�VR�Ћ�8�Q�J�E�P�у���^��]���������������U�졸8��$��SVu��8�H�1���8�J<�URP�A�Ѓ�����8�Q�J�E�P�ы�8�B�P�M�QV�ҡ�8�H�A�U�R�Ћ�8�Q�Jj j��E�h�*P�ы�8�B�@@�� j �M�Q�U�R�M��Ћ�8�Q�J���E�P���у���t/��8�B�u�HV�ы�8�B�P�M�Q�҃���^[��]á�8�P�E��RHjP�M��ҡ�8�P�E�M��RLj�j�PQ�M��ҡ�8�H�A�U�R�Ћ�8�Q�Jj j��E�h�*P�ы�8�B�@@��j �M�Q�U�R�M��Ћ�8�Q�J���E�P���у����3�����8�P�E��RHjP�M��ҡ�8�P�E�M��RLj�j�PQ�M��ҡ�8�H�u�QV�ҡ�8�H�A�U�VR�Ћ�8�Q�J�E�P�у���^[��]����������������U�졸8��$��SVu��8�H�1���8�J<�URP�A�Ѓ�����8�Q�J�E�P�ы�8�B�P�M�QV�ҡ�8�H�A�U�R�Ћ�8�Q�Jj j��E�h�*P�ы�8�B�@@�� j �M�Q�U�R�M��Ћ�8�Q�J���E�P���у���t/��8�B�u�HV�ы�8�B�P�M�Q�҃���^[��]á�8�P�E��RHjP�M��ҡ�8�P�E�M��RLj�j�PQ�M��ҡ�8�H�A�U�R�Ћ�8�Q�Jj j��E�h�*P�ы�8�B�@@��j �M�Q�U�R�M��Ћ�8�Q�J���E�P���у����3�����8�P�E��RHjP�M��ҡ�8�P�E�M��RLj�j�PQ�M��ҡ�8�H�A�U�R�Ћ�8�Q�Jj j��E�h�*P�ы�8�B�@@��j �M�Q�U�R�M��Ћ�8�Q�J���E�P���у����������8�P�E��RHjP�M��ҡ�8�P�E�M��RLj�j�PQ�M��ҋu�E�P���������8�Q�J�E�P�у���^[��]�������U�졸8��$��SVu��8�H�1���8�J<�URP�A�Ѓ�����8�Q�J�E�P�ы�8�B�P�M�QV�ҡ�8�H�A�U�R�Ћ�8�Q�Jj j��E�h�*P�ы�8�B�@@�� j �M�Q�U�R�M��Ћ�8�Q�J���E�P���у���t/��8�B�u�HV�ы�8�B�P�M�Q�҃���^[��]á�8�P�E��RHjP�M��ҡ�8�P�E�M��RLj�j�PQ�M��ҡ�8�H�A�U�R�Ћ�8�Q�Jj j��E�h�*P�ы�8�B�@@��j �M�Q�U�R�M��Ћ�8�Q�J���E�P���у����3�����8�P�E��RHjP�M��ҡ�8�P�E�M��RLj�j�PQ�M��ҡ�8�H�A�U�R�Ћ�8�Q�Jj j��E�h�*P�ы�8�B�@@��j �M�Q�U�R�M��Ћ�8�Q�J���E�P���у����������8�P�E��RHjP�M��ҡ�8�P�E�M��RLj�j�PQ�M���j h�*�M��b�����8�P�R@j �E�P�M�Q�M��҅���8�H�A�U�R���Ѓ���t/��8�Q�u�BV�Ћ�8�Q�J�E�P�у���^[��]Ë�8�M��B�PHjQ�M��ҡ�8�P�E�M��RLj�j�PQ�M��ҋu�E�P��������8�Q�J�E�P�у���^[��]���������������U���8�H<�A]����������������̡�8�H<�Q�����V��~ u>���t��8�Q<P�B�Ѓ��    W�~��t���:  W�  ���F    _^��������U���V�E�P���N�  ��P��������M����~  ��^��]��̃=�8 uK��8��t��8�Q<P�B�Ѓ���8    ��8��tV���~  V��  ����8    ^������������U���8��8�H�AS�U�V3�R�]��Ћ�8�Q�JSj��E�h�*P�ы�8�B<�P�M�Q�ҋ��8�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��xL �M�Q�U�R�M���L ����   W�}�}���   ��8���   �U��ATR�Ћ�����tB��8�Q�J�E�P���у��U�Rj�E�P��������8�Q�ȋBxW�Ѕ��E�t�E� ��t��8�Q�J�E�P����у���t��8�B�P�M�Q����҃��}� u"�E�P�M�Q�M���K ���;����E�_^[��]ËU��U�_�E�^[��]��������������U���DSV�u3�;�]�u_��8�H�A�U�R�Ћ�8�Q�JSj��E�h�*P�ы�8�B<�P�M�Q�ҋ��8�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]���J �M�Q�U�R�M��AK ���p  W�}��I �E����   ��8���   �U��ATR�Ћ�������   ��8�Q�J�E�P���ы�8�B���   ���M�Qj�U�R���Ћ�8�Q�J���E�P�ы�8�B�P�M�QV�ҡ�8�H�A�U�R�Ћ�8�Q�Bx��W�M��Ѕ��Et�E ��t��8�Q�J�E�P����у���t��8�B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*��8���   P�BH�Ћ�8�Q���ȋBxW�Ѕ�t"�M�Q�U�R�M���I ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M��CI �EP�M�Q�M�u��u�I ����   �u���E���tA��t<��uZ��8���   �M�PHQ�ҋ�8�Q���ȋBxV�Ѕ�u-�   ^��]Ë�8���   �E�JTP��VP�[�������uӍUR�E�P�M��I ��u�3�^��]����������V��~ u>���t��8�Q<P�B�Ѓ��    W�~��t����y  W�D  ���F    _^�������̋�� �*����������*���������̅�t��j�����̡�8�P��  ���8�P��(  ��U���8�P��   ��V�E�P�ҋuP���*y  �M��by  ��^��]� ��������̡�8�P��$  ��U���8�H��  ]��������������U���8�H���  ]�������������̡�8�H��  ��U���8�H���  ]��������������U���8�H��x  ]��������������U���8�H��|  ]��������������U���EV����*t	V��  ����^]� �������������̸   � �������̸   @� �������̸   � �������̸   � ��������U���8�H�QV�uV�҃���^]� �3�� �����������3�� �����������U����   h�   ��@���j P�TD �M�Eh�   ��@���R�M��MPQjǅ`���    ��  �� ��]���U����   V�u��u3�^��]�h�   ��@���j P��C �M�U�Eh�   �M���@���Q�U��U��@����ERPj��`���ǅD���PJ�E��N�E� �E� O�E�O�E��u�E��u�E�`%�D  �� ^��]�������������U���   SV�u(3ۅ��]�u��8�H�A�UR�Ѓ�^3�[��]Ë�8�Q�B<W�M3��Ѕ��'  �F ���E�tq�MQ�M���u  Wh�*�M��[���P�M���u  �u�Wj��U�R�E�P��\���Q�_?腉  ��P��x���R�y  ��P�E�P�y  ��P���MG ���E�t�E� �� t�M����� v  ��t��x��������u  ��t��\��������u  ��t�M̃����u  ��t��8�Q�J�E�P����у���t�M��u  �}� t"�U(�E$�M�R�UP�EQ�MRPQ����������U�R��D ����E$�M�UVP�Ej QRP�����������8�Q�J�EP�у���_^[��]���������������̋�`����������̋�`����������̋�`�����������U��V�u���t��8�QP��Ѓ��    ^]���������̡�8�H��@  hﾭ���Y����������U��E��t��8�QP��@  �Ѓ�]����������������U���8�H���  ]��������������U���8�H��  ]�������������̡�8�H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW�P ������u_^]Ã} tWj V�\@ ��_������F��8   ^]���U���8�ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW�2P ������u_^]�Wj V��? ��_������F��8   ^]�������������U���8�ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW�O ������u_^]�Wj V�f? ��_������F��8   ^]�������������U���8�ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW�2O ������u_^]�Wj V��> ��_������F��8   ^]�������������U���8�ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW�N ������u_^]�Wj V�f> ��_������F��8   ^]�������������U��M��t-�=�8 t�y���A�uP�O ��]á�8�P�Q�Ѓ�]��������U��M��t-�=�8 t�y���A�uP��N ��]á�8�P�Q�Ѓ�]��������U���8�H�U�R�Ѓ�]���������U���8�H�U�R�Ѓ�]���������U���8�ɋEt#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�nM ������u_^]�Wj V�"= ��_������F��8   ^]���������U���8�ɋEtL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËMQ������]�������U��E��w�   ��8��t�U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�L ������u_^]�Wj V�3< ��_������F��8   ^]����������U��E��w�   ��8��t,�} �U�IR�URPt���   �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW��K ������u_^]�Wj V�; ��_������F��8   ^]�������U���8�H�U�R�Ѓ�]���������U���8�H�U�R�Ѓ�]���������U���8�H�U�R�Ѓ�]���������U���8�H�U�R�Ѓ�]���������U���8�Hp�]���8�Hp�h   �҃�������������U��V�u���t��8�QpP�B�Ѓ��    ^]���������U���8�Pp�EP�EPQ�J�у�]� U���8�Pp�EP�EPQ�J�у�]� U���8�Pp�EP�EPQ�J�у�]� U���8�Pp�EPQ�J�у�]� ����U��E��8� ]��U���8�P8�EPQ�JD�у�]� ���̡�8�H8�Q<�����U���8�H8�A@V�u�R�Ѓ��    ^]�������������̡�8�H8�������U���8�H8�AV�u�R�Ѓ��    ^]��������������U���8�P8�EP�EP�EPQ�J�у�]� ������������U���8�P8�EP�EPQ�J�у�]� ��8�P8�BQ�Ѓ����������������U���8�P8�EPQ�J �у�]� ����U���8�P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U���8�P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U���8�P8�EP�EPQ�J(�у�]� U���8�P8�EP�EP�EPQ�J,�у�]� ������������U���8�P8�EP�EP�EPQ�J�у�]� ������������U���8�P8�EP�EP�EP�EP�EPQ�J�у�]� ����U���8�P8�EP�EPQ�J0�у�]� U���8�P8�EP�EP�EPQ�J4�у�]� ������������U���8�P8�EPQ�J8�у�]� ����U���8�H��x  ]��������������U���8�H��|  ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H�A,]�����������������U���8�H�QV�uV�ҡ�8�H�Q8V�҃���^]�����̡�8�H�Q<�����U���8�H�I@]����������������̡�8�H�QD����̡�8�H�QH�����U���8�H�AL]�����������������U���8�H�IP]�����������������U���8�H��<  ]��������������U���8�H��,  ]��������������U���8�H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡�8�H���   ���8�H���  ��U���8�H�U�ER�UP�ER�UP���   Rh�.  �Ѓ�]����������������U���8�H�A]�����������������U���8�H��\  ]��������������U���8�H�AT]�����������������U���8�H�AX]�����������������U���8�H�A\]����������������̡�8�H�Q`����̡�8�H�Qd����̡�8�H�Qh�����U���8�H�Al]�����������������U���8�H�Ap]�����������������U���8�H�At]�����������������U���8�H��D  ]��������������U���8�H��  ]��������������U���8�H�Ix]�����������������U���8�H��@  ]��������������U��V�u����e  ��8�H�U�A|VR�Ѓ���^]���������U���8�H���   ]��������������U���8�H��h  ]��������������U���8�H��d  ]��������������U���8�H���  ]�������������̡�8�H���   ��U���8�H��l  ]��������������U���8�H��   ]��������������U���8�H��  ]��������������U��V�u���r�  ��8�H���   V�҃���^]���������̡�8�H��`  ��U���8�H��  ]��������������U���8�H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U���8�H���  ]��������������U��U�E��8�H�E���   R���\$�E�$P�у�]�U���8�H���   ]��������������U���8�H���   ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H���   ]��������������U���8�H���   ]��������������U���8�H���   ]��������������U���8�H���   ]��������������U���8�H���   ]��������������U���8�H���   ]��������������U���8�P���E�P�E�P�E�PQ���   �у����#E���]����������������U���8�P���E�P�E�P�E�PQ���   �у����#E���]����������������U���8�P���E�P�E�P�E�PQ���   �у����#E���]����������������U���8�H��8  ]��������������U��V�u(V�u$�E�@��8�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@��8�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U���8�P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U���8�P0�EP�EP�EP�EPQ���   �у�]� ����̡�8�P0���   Q�Ѓ�������������U���8�P0�EP�EPQ���   �у�]� �������������U���8�P0�EP�EP�EP�EPQ���   �у�]� ����̡�8�P0���   Q�Ѓ������������̡�8�H0���   ��U���8�H0���   V�u�R�Ѓ��    ^]�����������U���8�H��H  ]��������������U���8�H��T  ]�������������̡�8�H��p  ���8�H���  ��U���8�H���  ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H�U�E��X  ��VR�UPR�E�P�ыu�    �F    ��8���   �Qj PV�ҡ�8���   ��U�R�Ѓ� ��^��]��������U���$Vj hLGOg�M���  P�E�hicMCP�k������M���  ��8���   �JT�E�P�у���u(�u��芺  ��8���   ��M�Q�҃���^��]á�8���   �AT�U�R�Ћu��P��芺  ��8���   �
�E�P�у���^��]�������������U���8�H��  ]��������������U���8�H��\  ]��������������U���8�H�U��t  ��V�uVR�E�P�у����^  �M���]  ��^��]�����U���8�H�U���  ��VWR�E�P�ы�8�u���B�HV�ы�8�B�HVW�ы�8�B�P�M�Q�҃�_��^��]����������������U���8�H�U���  ��VWR�E�P�ы�8�u���B�HV�ы�8�B�HVW�ы�8�B�P�M�Q�҃�_��^��]����������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H�U�E��VWj R�UP�ERP��t  �U�R�Ћ�8�Q�u���BV�Ћ�8�Q�BVW�Ћ�8�Q�J�E�P�у�(_��^��]��U���8�H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    ��8���   j P�BV�Ћ�8���   �
�E�P�у�$��^��]���U���8�H��8  ]��������������U���  �  3ŉE��M�EPQ������h   R�b ����|	=�  |#���8�H��0  h�*hF  �҃��E� ��8�H��4  ������Rh,+�ЋM�3̓��" ��]�������U���8�H��  ��V�U�WR�Ћ�8�Q�u���BV�Ћ�8�Q�BVW�Ћ�8�Q�J�E�P�у�_��^��]����U���8�H��  ��V�U�WR�Ћ�8�Q�u���BV�Ћ�8�Q�BVW�Ћ�8�Q�J�E�P�у�_��^��]����U���8�H��p  ��$�҅�trh���M��ɵ  ��8�P�E�R4Ph���M��ҡ�8�P�E�R4Ph���M���j �E�P�M�hicMCQ������8���   ��M�Q�҃��M�褵  ��]�U���8�H��p  ��$V�҅�u��8�H�u�QV�҃���^��]�Wh!���M���  ��8�P�E�R4Ph!���M���j �E�P�M�hicMCQ������8���   �QHP�ҋu����8�H�QV�ҡ�8�H�QVW�ҡ�8���   ��U�R�Ѓ�$�M��ݴ  _��^��]������U���8�H��p  ��$V�҅�u��8�H�u�QV�҃���^��]�Wh����M��L�  ��8�P�E�R4Ph����M���j �E�P�M�hicMCQ������8���   �QHP�ҋu����8�H�QV�ҡ�8�H�QVW�ҡ�8���   ��U�R�Ѓ�$�M���  _��^��]������U���8�H��p  ��$�҅�u��]�Vh#���M�蔳  ��8�P�E�R4Ph#���M���j �E�P�M�hicMCQ�������8���   �Q8P�ҋ��8���   ��U�R�Ѓ��M��u�  ��^��]���������������U���8�H��p  ��$�҅�u��]�Vhs���M����  ��8�P�E�R4Phs���M���j �E�P�M�hicMCQ�W�����8���   �Q8P�ҋ��8���   ��U�R�Ѓ��M��ղ  ��^��]���������������U���8�H���  ]��������������U���8�H��@  ]��������������U���8�H���  ]��������������U��V�u���t��8�QP��D  �Ѓ��    ^]������U���8�H��H  ]��������������U���8�H��L  ]��������������U���8�H��P  ]��������������U���8�H��T  ]��������������U���8�H��X  ]��������������U���8�H��\  ]�������������̡�8�H��d  ��U���8�H��h  ]��������������U���8�H��l  ]�������������̡�8�H���  ��U���8�H�U���  ��VR�E�P�ыu��P���ð  �M��۰  ��^��]�����U���8�H���  ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H���  ]��������������U���8�H��$  ]��������������U���8�H��(  ]��������������U���8�H��,  ]�������������̡�8�H��0  ���8�H��<  ��U���8�H���  ]�������������̡�8�H���  ��U���8�H���  ]������������������������������U���8�H��  ]�������������̡�8�H��P  ���8���   ���   ��Q��Y��������U���8�H�A�U��� R�Ћ�8�Q�Jj j��E�h0+P�ыUR�E�P�M�Q�-�����8�B�P�M�Q�ҡ�8�H�A�U�R�Ћ�8�Q�J�E�P�у�,��]�̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������U���   V���O  �����   �ESP�M��8P  ��8�Q�J�E�P�ы�8�B�Pj j��M�h�*Q�҃��E�P�M���O  j j��M�Q�U�R��d���P�c  ��P�M�Q�S  ��P�U�R�S  ���P�o! ���M����1P  �M��)P  ��d����P  �M��P  ��8�H�A�U�R�Ѓ��M���O  ��[t	V� ����^��]� ���U��EVP����) �����^]� �����Q�J Y���������U��E�M�U�H4�M�P �U��M�@PJ�@8�N�@<`%�@@ �@D�u�@H�u�@L O�@P�u�@l��@X�u�@\��@`�u�@d��@TO�@h �@p��@t�u�P0�H(�@,    ]��������������U���   h�   ��`���j P�t �M�U�Ej Q�MRPQ��`���R�����E �Uh�   ��`���Q�E��ERPj�������8��]��������������̋�`����������̋�` ����������̋�`@����������̋�`����������̋�`8����������̋�`,�����������h�8PhD ��0 ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d��������]� ���������U��h�8jhD ��/ ����t
�@��t]��3�]��������Vh�8j\hD ���/ ����t�@\��tV�Ѓ���^�����Vh�8j`hD ���/ ����t�@`��tV�Ѓ�^�������U��Vh�8jdhD ���Y/ ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh�8jhhD ���/ ����t�@h��t
�MQV�Ѓ�^]� ������������Vh�8jlhD ����. ����t�@l��tV�Ѓ�^�������U��Vh�8h�   hD ���. ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�8h�   hD ���V. ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�8jphD ���	. ����t�@p��t�MQV�Ѓ�^]� ��8^]� ��U��Vh�8jxhD ����- ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh�8j|hD ���- ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh�8j|hD ���I- ����t�@|��t�MVQ�Ѓ������^]� �   ^]� ����������̋���������������h�8jhD ��, ����t	�@��t��3��������������U��V�u�> t+h�8jhD �, ����t�@��tV�Ѓ��    ^]�������U��VW�}����t0h�8jhD �q, ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh�8jhD ���), ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh�8jhD ����+ ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh�8j hD ���+ ����t�@ ��tV�Ѓ�^�3�^���Vh�8j$hD ���|+ ����t�@$��tV�Ѓ�^�3�^���U��Vh�8j(hD ���I+ ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh�8j,hD ����* ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh�8j(hD ���* ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh�8j4hD ���l* ����t�@4��tV�Ѓ�^�3�^���U��Vh�8j8hD ���9* ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh�8j<hD ����) ����t�@<��t
�MQV�Ѓ�^]� ������������Vh�8jDhD ���) ����t�@D��tV�Ѓ�^�3�^���U��Vh�8jHhD ���y) ����t�M�PHQV�҃�^]� U��Vh�8jLhD ���I) ����u^]� �M�PLQV�҃�^]� �����������U��Vh�8jPhD ���	) ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh�8jThD ����( ����u^Ë@TV�Ѓ�^���������U��Vh�8jXhD ���( ����t�M�PXQV�҃�^]� U��Vh�8h�   hD ���f( ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh�8h�   hD ���( ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh�8h�   hD ����' ����u^]� �M���   QV�҃�^]� �����U��Vh�8h�   hD ���' ����u^]� �M���   QV�҃�^]� �����U��Vh�8h�   hD ���F' ����u^]� �M���   QV�҃�^]� �����U��Vh�8h�   hD ���' ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh�8h�   hD ��& ����u��8�H�u�QV�҃���^��]ËM���   WQ�U�R�Ћ�8�Q�u���BV�Ћ�8�Q�BVW�Ћ�8�Q�J�E�P�у�_��^��]��U��Vh�8h�   hD ���6& ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�8h�   hD ����% ����t���   ��t�MQ����^]� 3�^]� �U��Vh�8h�   hD ���% ����t���   ��t�MQ����^]� 3�^]� �U��Vh�8h�   hD ���f% ����t���   ��t�MQ����^]� 3�^]� �Vh�8h�   hD ���)% ����t���   ��t��^��3�^����������������U��Vh�8h�   hD ����$ ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�8h�   hD ���$ ����t���   ��t�MQ����^]� ��������U��Vh�8h�   hD ���V$ ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vh�8h�   hD ���	$ ����t���   ��t��^��3�^����������������VW��3����$    �h�8jphD �# ����t�@p��t	VW�Ѓ����8�8 t����_��^�����U��SW��3�V��    h�8jphD �o# ����t�@p��t	WS�Ѓ����8�8 tsh�8jphD �=# ����t�@p��t�MWQ�Ѓ������8h�8jphD �# ����t�@p��t	WS�Ѓ����8V���7�����t���[����E��^t�8��~=h�8jphD �" ����t�@p��t	WS�Ѓ����8�8 u_�   []� _3�[]� ��������U��Vh�8j\hD ���i" ����t3�@\��t,V��h�8jxhD �G" ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh�8j\hD ���	" ����t3�@\��t,V��h�8jdhD ��! ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh�8j\hD ���! ����tG�@\��t@V�ЋEh�8jdhD �E��E�    �E�    �p! ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh�8j\hD ���)! ����t\�@\��tUV��h�8jdhD �! ����t�@d��t
�MQV�Ѓ�h�8jhhD ��  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh�8j\hD ���  ������   �@\��t~V��h�8jdhD �s  ����t�@d��t
�MQV�Ѓ�h�8jhhD �J  ����t�@h��t
�URV�Ѓ�h�8jhhD �!  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh�8jthD ���� ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h�8j`hD � ����t(�@`��t!�M�Q�Ѓ���^��]� �uh�8���_�����^��]� ������U���Vh�8h�   hD ���S ����tR���   ��tH�MQ�U�R���ЋuP������h�8j`hD � ����t<�@`��t5�M�Q�Ѓ���^��]� �u�U�R���E�    �E�    �E�    ������^��]� ��������������U�����E��������u
���@+]��0'������u
���8+]�]�D ����U��V�u�������E���P�V�H�N�P�V�H�N�P�V��^]���������U��V�u������E� �^�@�^8�@���^X^]����������U���V�u��菗���E�W �]��E�| �E��VX�������^@���^P�^8^��]�U���V�u���O����E� �]��E�< �E��V�������^H���^(�^X^��]�U���V�u�������E�� �]��E�� �E��V�����V0���^ �^8^��]���U�������e�5H+�U��$� �m��H+�������E���$������Az
���.���]��؋�]��������������U���`�E� ���$�P��V�ɉM�H�]ЉU�P��W�`�}�M��H�]؉U�P�@���u�M��]��U���$�B����]��u��G�$�1����]��u��G�$� ����]ȍu���$�����]��u��G�$������]��u��G�$������E�����_�E�^�����������E����E������E�����������A�Eu�E���E��X�E��X��]ËM�U��M��P�U�H�M��P�U��H�P��]�������������U�����V�u�V�VW�}��G����������f �U��P+������Au>�����W��������z�@+_����^�^^��]��8+_����^�^^��]�����_���?���$z	�m�������d�����$����G�u��� �^��_�^��^��]���������������U���PV�u�FP�M�Q�.���FH�U����FP�]��FX�U���������� �U��P+^������A��   �����U��E����E��E���������������Az�����)�0'������u
����$������e �E����������U�����z1�@+���������D  �E���H+���E���X�X��]��8+��������A�  �E���H+���E���X�X��]�����]����}����$z	��������������$�U�����������Au�H+�]�����E��u��| �]��E��� �]��E�� �E��M��E������������M�����������Az�����$�0'������u
����$����= ���������]�����z�E���-H+�E��E���X�X��]ËE���E��E���X�X��]ËE���E���X�X��]����U�����   V���u�����Dz%�V����Dz�^����Dz�u���(�����^��]�����U�� �]��E��� ݝx����F�U��� �]��E�� ݝp����F�U��� �]��E�� �E����  �$���E�u���E��E�P�ɍM�݅x���Q�ˍU�R�E���P�E��������������]������������]�݅p��������]������]������]��E����]������������]��������������]����]����U��U��]�蕑����^��]��E��M���Q݅x����U���R�E��E���P�ˍM�Q�U��������]�݅p������E����������]������E������]��E��]������]��������]��������]������������]��  ���U��E�R�ɍE��E�P���M���Q�U�R�U������]��E���݅x��������]�݅p��������]������]������������]��E����������]������]������������]����  �E��E���P݅p����M���Q�E�U���R�ˍE�P�U�݅x��������E��������]������]��E����������]������������]��������]������������]����]��E����]����  �E�M���Q�E��U���R݅p����E���P�ʍM��E�Q�����������]������������]���݅x��������]������������]������������]��������]������]������]��E��   ���U��E�R�ɍE��E�P���M���Q�U�R�]�݅p������E��������]����]���݅x��������]������������]������]��������������]������E����������]��������]������������u�]�����U��U��]��ʎ����^��]ÍI ��"���=�+�����������U���xV�uW�   �}��E��P�M�Q�>(����H�U��P�M��H�U��P�@�M��M��U�Q�U�R�E��(����P�M��H�U��P�M��H�UċP�EЉM�P�M�Q�U���'���E���E��H�UЋP�MԋH�U؋P�@�E�U��E������M�����$��������u������0'������u
����$��� �}�u��EȍM��e�VQ��E��e��^�E��e��^�H'������H�N�P�V�H�N�P�V�@�F�������Dz,�V����Dz"�V����Dz����������^�^�_^��]�_��^��]�����U���0V�uW��螌����}�������Dz�W����Dz
�W����D{�E��������Dz
_�؋�^��]���$�U��T �]��E�� �]��E�WP�l&��� �E������@���@�����X+�������������E������]������]������������]��������������������������]��E����]����E������]��E��^�E��^ �E��^(�E������]��������������]����E�����_�]����E��^0�E��^8�E��^@���������������^H���^P�^X^��]��������������U��E�A    �]� �������������U��Q���i�� %������E���E�}�h+�5`+��]�U��Q���i�� %������E���E�}�h+�5`+���%�$��]���������U���V��~ ��   �`+��X+������؍Ai�� %����ȅɉM��E�}�h+��Hi�� ���������U��х҉U��E�}�h+�������U����������U�������t���������D{��ډ������� �x+�u��H� �E����F   �^^�M��p+��$��]��F�F    �p+^��$��]�����������U���V��~ ��   �`+��X+������؍Ai�� %����ȅɉM��E�}�h+��Hi�� ���������U��х҉U��E�}�h+�������U����������U�������t���������D{��ډ������� �x+�u��H� �E����F   �^^�M���+��]��F�F    ��+^��]�������U��E�M�@�I�����A�H����� ���@�����H�E�������A�����X�i�X]�������U��E� �@�@����������Au��������������Au����������������z��������������z����������������   ����������'������Au�E������������X�X]�������������Dz
���������5��������Dz�������������X+��������������H'�������5�+��������z��$�E����X�X]ËE�����������P�P�]�U����E� �@�U��@�U���'��������Au�E������������X�X��]�����������Dz������+���U��$�� �E����������E����E������������������������������ �����wE�$�̙�����ʋE��������X�X��]��������������ۋE��������X�X��]����������������U��M�A��A��������������������������Dz�E���P�P�]ËU�؋E�� �B�`�B�`������I���I����������I���I� �����@�@�E���������j�X�j�X]�������̡�8�H���   ��U���8�H���   V�u�R�Ѓ��    ^]����������̡�8�H���   ��U���8�H���   V�u�R�Ѓ��    ^]����������̡�8�P���   Q��Y��������������U��� ��8SV��H�QPWV�u�����}�W�W3����;��W(�W �E��_��$�_0����������_�_��$�������_���_ �_(~w��u���8�H�QLSV�ҋ����<t<uL�F(�E��f@P���]��F0�fH�]��F8�fP�]��y����F@�M��F(Q���]��F0�FH�]��F8�FP�]��S�����;]�|���_^[��]� U���8�P�EPQ���   �у�]� �U���8�P�EP�EP�EP�EP�EP�EPQ���   �у�]� �������������U���8�P�EP�EP�EP�EP�EP�EPQ���   �у�]� �������������U���8�P�EP�EP�EP�EPQ���   �у�]� �����U���8�P�EP�EP�EP�EPQ��  �у�]� �����U���8�P�EP�EP�EP�EPQ���  �у�]� �����U���8�P�EP�EPQ���   �у�]� �������������U��V�uW�����o�  ��8�H���   VW�҃�_��^]� ��U���8�P�EPQ���   �у�]� �U���8�P�EPQ��  �у�]� ̡�8�P��0  Q�Ѓ�������������U���8�P�EP�EPQ��t  �у�]� �������������U���8�H�U���  j R�Ѓ�]���U���8�H���  V�u�R�Ѓ��    ^]�����������U���8�H���   ]��������������U���8�H���   V�u�R�Ѓ��    ^]�����������U��� ���83��U�Q�U�Q�]�Q�M��M��P�E�PQ�E�P�EPPP�EP�EP�EP�EPQ��d  �у�8��]��������������U��U��tA���    t8��  �M;A}*V�1�0^t	�E�    �	��  �t	�E�    ]����U���8�H��P  ]��������������U���8�H��T  ]��������������U���8�H��X  ]�������������̋��     ��������V����t��8�QP��<  �Ѓ��    ^�����������U����t��8�Q�M���  Q�MQP�҃�]� ������U����t��8�Q�M���  Q�MQP�҃�]� ������U���8��S3�V��W�};���~D�^<�^8�^@�^H�FL   �^P�^T��   �U�R���
  P�N�o&  �M��7#  ����  �F�E�P���  ��N�P�V�H�N�P�V��8�H@�Q,W�ҋ���;�tG��8�P���   Sh6  ���ЉFP��8�Q���   Sh5  ����_�FT^[��]� �F   _^[��]� ���̋��@    � d   �V����t��8�QP��<  �Ѓ��    ^�����������U��V����t��8�QP��<  �Ѓ��    ��8�Q�E�MP�EQ��8  P��3҃����^��]� ��������̡�8�HL���   ��U���8�H@�AV�u�R�Ѓ��    ^]�������������̡�8�HL�������U���8�H@�AV�u�R�Ѓ��    ^]�������������̡�8�PL���   Q�Ѓ�������������U���8�PL�EP�EPQ���   �у�]� �������������U���8V��HL���   V�҃���u��8�U�HL���   j RV�Ѓ�^]� ��8���   �ȋBP�Ћ�8���   �MP�BH��^]� �����̡�8�PL��(  Q�Ѓ�������������U���8�PL�EP�EPQ��,  �у�]� ������������̡�8�HL�Q�����U���8�H@�AV�u�R�Ѓ��    ^]��������������U���8�PL�E�R��VPQ�M�Q�ҋu��P���%|  �M��=|  ��^��]� ����U���8�PL�EPQ���   �у�]� �U���8�PL�EP�EPQ�J�у�]� ��8�PL�BQ�Ѓ���������������̡�8�PL�BQ�Ѓ���������������̡�8�PL�BQ�Ѓ����������������U���8�PL�EP�EP�EPQ�J �у�]� ������������U���8�PL�EPQ��4  �у�]� �U���8�PL�EP�EP�EPQ�J$�у�]� ������������U���8�PL�EP�EP�EP�EPQ�J(�у�]� �������̡�8�PL�B,Q�Ѓ���������������̡�8�PL�B0Q�Ѓ����������������U���8�PL�EP�EPQ��  �у�]� ������������̡�8�PL���   Q�Ѓ�������������U���8�PL�E��  ��VPQ�M�Q�ҋu��P���z  �M��z  ��^��]� ̡�8�PL�B4Q�Ѓ���������������̡�8�PL�B8j Q�Ѓ��������������U���8�PL���   ]��������������U���8�PL���   ]��������������U���8�PL���   ]��������������U���8�PL���   ]��������������U���8�PL���   ]��������������U���8�PL���   ]��������������U���8�PL���   ]��������������U���8�PL���   ]��������������U���8�PL���   ]��������������U���8�PL�EPQ�J<�у�]� ���̡�8�PL�BQ��Y�U���8�PL�EP�EPQ�J@�у�]� U���8�PL�Ej PQ�JD�у�]� ��U���8�PL�Ej PQ�JH�у�]� ��U���8�PL�EjPQ�JD�у�]� ��U���8�PL�EjPQ�JH�у�]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}������W�M�Q�U�R����A  ���M����W�����t��8���   ��U�R�Ѓ�_^3�[��]Ë�8���   �J8�E�P�ы�8�����   ��M�Q�҃�_��^[��]��������������U���$3�V�E��E�E��P�M��E�   �E�   �E��  �>���j�M�Q�U�R���MA  �M�������8���   ��U�R�Ѓ�^��]�����������U���$��8�UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}�����j�E�P�M�Q����@  �M��!�����8���   ��M�Q�҃�_^��]� ��U���$��8�UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��:���j�E�P�M�Q���I@  �M�������8���   ��M�Q�҃�_^��]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}������W�M�Q�U�R����?  ���M����7�����t+�u���9  ��8���   ��U�R�Ѓ�_��^[��]� ��8���   �JL�E�P�ыu��P���  ��8���   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}�����W�M�Q�U�R���?  ���M����w�����t+�u���y  ��8���   ��U�R�Ѓ�_��^[��]� ��8���   �JL�E�P�ыu��P����  ��8���   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��T���W�M�Q�U�R���D>  ���M�������_^��[t��8���   ��U�R�������]Ë�8���   �J<�E�P���]���8���   ��M�Q���E�����]���������������U���$SVW3��E��P�M��}܉}��E��  �}��}�����W�M�Q�U�R���=  ���M���������t��8���   ��U�R�Ѓ�_^3�[��]Ë�8���   �J8�E�P�ы�8�����   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}������W�M�Q�U�R����<  ���M����W�����t-��u��8����   ���^�U�R�Ѓ�_��^[��]� ��8���   �JP�E�P�ы�u�H��P�@�N��8�V���   �
�F�E�P�у�_��^[��]� �����̡�8�PL���   Q��Y��������������U���8�PL�E���   ��jPQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���8�PL�E���   ��j PQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���$SVW3��E��P�M��}܉}��E��  �}��}��d���W�M�Q�U�R���T;  ���M����������t-��u��8����   ���^�U�R�Ѓ�_��^[��]� ��8���   �JP�E�P�ы�u�H��P�@�N��8�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}�����W�M�Q�U�R���:  ���M����������t-��u��8����   ���^�U�R�Ѓ�_��^[��]� ��8���   �JP�E�P�ы�u�H��P�@�N��8�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}������W�M�Q�U�R���9  ���M����'�����t-��u��8����   ���^�U�R�Ѓ�_��^[��]� ��8���   �JP�E�P�ы�u�H��P�@�N��8�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}������W�M�Q�U�R����8  ���M����W�����t��8���   ��U�R�Ѓ�_^3�[��]Ë�8���   �J8�E�P�ы�8�����   ��M�Q�҃�_��^[��]��������������U����E3�V�]�E��E��E��P�M�E�   �E��  �?���j�M�Q�UR���N8  �M������8���   ��U�R�Ѓ�^��]� ���������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E������j�U�R�E�P����7  �M��6�����8���   �
�E�P�у�^��]� ��������U���$��8�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��J���j�E�P�M�Q���Y7  �M�������8���   ��M�Q�҃�_^��]� ��U���$��8�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}������j�E�P�M�Q����6  �M��1�����8���   ��M�Q�҃�_^��]� ��U���$��8�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��J���j�E�P�M�Q���Y6  �M�������8���   ��M�Q�҃�_^��]� ��U���$��8�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}������j�E�P�M�Q����5  �M��1�����8���   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��_���j�U�R�E�P���n5  �M��������8���   �
�E�P�у�^��]� ��������U���$SVW3��E��P�M��}܉}��E��  �}��}������W�M�Q�U�R����4  ���M����W�����t-��u��8����   ���^�U�R�Ѓ�_��^[��]� ��8���   �JP�E�P�ы�u�H��P�@�N��8�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��$���W�M�Q�U�R���4  ���M���������t��8���   ��U�R�Ѓ�_^3�[��]Ë�8���   �J8�E�P�ы�8�����   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��t���W�M�Q�U�R���d3  ���M����׿����t��8���   ��U�R�Ѓ�_^3�[��]Ë�8���   �J8�E�P�ы�8�����   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ����U���$��8�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}�����j�E�P�M�Q���2  �M�������8���   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E�����j�U�R�E�P���.2  �M�膾����8���   �
�E�P�у�^��]� ��������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E�����j�U�R�E�P���1  �M�������8���   �
�E�P�у�^��]� ��������U���8�H���   ]��������������U���8�H���   ]�������������̡�8�H���   ���8�H���   ��U���8�H���   V�u�R�Ѓ��    ^]�����������U���8�H���   ]��������������U���8�HL�QV�ҋ���u^]á�8�H�U�ER�UP���  RV�Ѓ���u��8�Q@�BV�Ѓ�3���^]����������U���8�H�U�E���  R�U�� P�ERP�у�]������U���8�H���   ]��������������U���8�H�U �ER�UP�ER�UP�ER�UP���   R�Ѓ�]������������̡�8�PL�BLQ�Ѓ���������������̡�8�PL�BPQ�Ѓ����������������U���8�PL�EP�EPQ�JT�у�]� U���8�PL�EPQ��  �у�]� �U���8�PL�EPQ���   �у�]� ̡�8�PL�BXQ�Ѓ����������������U���8�PL�EP�EP�EPQ�J\�у�]� ������������U���4��8SV��HL�QW�ҋ�3�;��}��x  �M��d  ��8�E�EԋE�]Љ]؉]܉]�]��}̋Q�R0Ph]  �M��ҡ�8���   �BSSW���Ѕ���   ��8�QL�BW�Ћ���;���   ��    ��8���   �B(���ЍM�Qh�   ���u�躠��������   �M�;���   ��8���   ���   S��;�tm��8���   �ȋB<V�Ћ�8���   ���   �E�P�у�;�t��8�B@�HV�у�;����\����}��M�葴���M��Ic  ��_^[��]� �}���8�B@�HW�ы�8���   ���   �M�Q�҃��M��I����M��c  _^3�[��]� �����̡�8�PL�B`Q�Ѓ���������������̡�8�PL�BdQ�Ѓ����������������U���8�PL�EPQ�Jh�у�]� ���̡�8�PL��D  Q�Ѓ������������̡�8�PL�BlQ�Ѓ����������������U���8�PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U$�EV�Ehp�hP�h0�h �R�Q�U R�UR�UR�U���A�$�5�8�vLRP���   Q�Ѓ�4^]�  ������̡�8�PL���   Q�Ѓ�������������U���8�PL�EP�EP�EPQ��   �у�]� ���������U���8�PL��H  ]�������������̡�8�PL��L  ��U���8�PL��P  ]��������������U���8�PL��T  ]��������������U���8�PL�EP�EP�EP�EP�EPQ���   �у�]� �U���8�PL�EP�EP�EPQ���   �у�]� ���������U���8�PL�EP�EP�EP�EPQ��   �у�]� �����U���8�HL���   ]��������������U���8�HL���   ]��������������U���8�HL���   ]�������������̡�8�HL��  ���8�HL��@  ��h9Ph^� ���  ���������������U��Vh9j\h^� ����  ����t�@\��t
�MQV�Ѓ�^]� ������������U��� ��8V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ};��E�t`;�t\��8�QLjP���   ���ЋM��U�Rh=���M�}�裛������8���   ���   �U�R�Ѓ��M��u��ܯ����_^��]Ë�8���   ���   �E�P�у��M��u�讯��_�   ^��]����U��� ��8V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ};��E�t`;�t\��8�QLjP���   ���ЋM��U�Rh<���M�}��Ӛ������8���   ���   �U�R�Ѓ��M��u�������_^��]Ë�8���   ���   �E�P�у��M��u��ޮ��_�   ^��]���̡�8V�񋈈   ���   V�҃��    ^���������������U���8�P�EP�EP�EPQ�J�у�]� �����������̡�8V��H�QV�ҡ�8�H$�QDV�҃���^�����������U���8V��H�QV�ҡ�8�H$�QDV�ҡ�8�U�H$�AdRV�Ѓ���^]� ��U���8V��H�QV�ҡ�8�H$�QDV�ҡ�8�U�H$�ARV�Ѓ���^]� ��U���8V��H�QV�ҡ�8�H$�QDV�ҡ�8�H$�U�ALVR�Ѓ���^]� �̡�8V��H$�QHV�ҡ�8�H�QV�҃�^�������������U���8�P$�EPQ�JL�у�]� ����U���8�P$�R]�����������������U���8�P$�Rl]����������������̡�8�P$�Bp����̡�8�P$�BQ�Ѓ����������������U���8�P$��VWQ�J�E�P�ы�8�u���B�HV�ы�8�B�HVW�ы�8�B�P�M�Q�҃�_��^��]� ���U���8�P$�EPQ�J�у�]� ����U���8�P$��VWQ�J �E�P�ы�8�u���B�HV�ы�8�B$�HDV�ы�8�B$�HLVW�ы�8�B$�PH�M�Q�ҡ�8�H�A�U�R�Ѓ� _��^��]� ���U���8�P$��VWQ�J$�E�P�ы�8�u���B�HV�ы�8�B$�HDV�ы�8�B$�HLVW�ы�8�B$�PH�M�Q�ҡ�8�H�A�U�R�Ѓ� _��^��]� ���U���V�uV�E�P�l������e�����8�Q$�JH�E�P�ы�8�B�P�M�Q�҃���^��]� ����̡�8�P$�B(Q��Yá�8�P$�BhQ��Y�U���8�P$�EPQ�J,�у�]� ����U���8�P$�EPQ�J0�у�]� ����U���8�P$�EPQ�J4�у�]� ����U���8�P$�EPQ�J8�у�]� ����U���8�UV��H$�ALVR�Ѓ���^]� ��������������U���8�H�QV�uV�ҡ�8�H$�QDV�ҡ�8�H$�U�ALVR�Ћ�8�E�Q$�J@PV�у���^]�U���8�UV��H$�A@RV�Ѓ���^]� ��������������U���8�P$�EPQ�J<�у�]� ����U���8�P$�EPQ�J<�у������]� �������������U���8�P$�EP�EPQ�JP�у�]� U���8�P$�EPQ�JT�у�]� ���̡�8�H$�QX�����U���8�H$�A\]�����������������U���8�P$�EP�EP�EPQ�J`�у�]� �����������̡�8�H(�������U���8�H(�AV�u�R�Ѓ��    ^]��������������U���8�P(�R]����������������̡�8�P(�B�����U���8�P(�R]�����������������U���8�P(�R]�����������������U���8�P(�R ]�����������������U���8�P(�E�RjP�EP��]� ��U���8�P(�E�R$P�EP�EP��]� ��8�P(�B(����̡�8�P(�B,����̡�8�P(�B0�����U���8�P(�R4]�����������������U���8�P(�RX]�����������������U���8�P(�R\]�����������������U���8�P(�R`]�����������������U���8�P(�Rd]�����������������U���8�P(�Rh]�����������������U���8�P(�Rx]�����������������U���8�P(�Rl]�����������������U���8�P(�Rt]�����������������U���8�P(�Rp]�����������������U���8�P(�BpVW�}W���Ѕ�t:��8�Q(�Rp�GP���҅�t"��8�P(�Bp��W���Ѕ�t_�   ^]� _3�^]� ��U���8�P(�BtVW�}W���Ѕ�t:��8�Q(�Rt�GP���҅�t"��8�P(�Bt��W���Ѕ�t_�   ^]� _3�^]� ��U��VW�}W���0�����t8�GP���!�����t)�OQ��������t��$W��������t_�   ^]� _3�^]� ������������U��VW�}W���0�����t8�GP���!�����t)�O0Q��������t��HW��������t_�   ^]� _3�^]� ������������U�����8�E�    �E�    �P(�RhV�E�P���҅���   �E���uG��8�H�A�U�R�Ћ�8�Q�E�RP�M�Q�ҡ�8�H�A�U�R�Ѓ��   ^��]� ��8�Qh�+h`  P���   �Ћ�8�����E��Q(u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P�f�����3�^��]� �M��U�j ���Q�MR�����E�P�<������   ^��]� �������������U���8��V��H�A�U�R�Ѓ��M�Q��������^u��8�B�P�M�Q�҃�3���]� ��8�H$�E�I�U�RP�ы�8�B�P�M�Q�҃��   ��]� �U��Q��8�P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U���8�P(�R8]�����������������U���8�P(�R<]�����������������U���8�P(�R@]�����������������U���8�P(�RD]�����������������U���8�P(�RH]�����������������U���8�P(�E�R|P�EP��]� ����U���8�P(�RL]�����������������U���8�E�P(�BT���$��]� ���U���8�E�P(�BPQ�$��]� ����̡�8�H(�Q�����U���8�H(�AV�u�R�Ѓ��    ^]��������������U���8�P(���   ]��������������U���8�H(�A]����������������̡�8�H,�Q,����̡�8�P,�B4�����U���8�H,�A0V�u�R�Ѓ��    ^]�������������̡�8�P,�B8�����U���8�P,�R<��VW�E�P�ҋu����8�H�QV�ҡ�8�H$�QDV�ҡ�8�H$�QLVW�ҡ�8�H$�AH�U�R�Ћ�8�Q�J�E�P�у�_��^��]� �������U���8�P,�E�R@��VWP�E�P�ҋu����8�H�QV�ҡ�8�H�QVW�ҡ�8�H�A�U�R�Ѓ�_��^��]� ��̡�8�H,�j j �҃��������������U���8�P,�EP�EPQ�J�у�]� U���8�H,�AV�u�R�Ѓ��    ^]�������������̡�8�P,�B����̡�8�P,�B����̡�8�P,�B����̡�8�P,�B ����̡�8�P,�B$����̡�8�P,�B(�����U���8�P,�R]�����������������U���8�P,�R��VW�E�P�ҋu����8�H�QV�ҡ�8�H$�QDV�ҡ�8�H$�QLVW�ҡ�8�H$�AH�U�R�Ћ�8�Q�J�E�P�у�_��^��]� �������U���8�H��D  ]��������������U���8�H��H  ]��������������U���8�H��L  ]��������������U���8�H�I]�����������������U���8�H�A]�����������������U���8�H�I]�����������������U���8�H�A]�����������������U���8�H�I]�����������������U���8�H���  ]��������������U���8�H�A]�����������������U���V�u�E�P���������8�Q$�J�E�P�у���u-��8�B$�PH�M�Q�ҡ�8�H�A�U�R�Ѓ�3�^��]Ë�8�Q�J�E�jP�у���u=�U�R��������u-��8�H$�AH�U�R�Ћ�8�Q�J�E�P�у�3�^��]Ë�8�B�HjV�у���u��8�B�HV�у����I�����8�Q$�JH�E�P�ы�8�B�P�M�Q�҃��   ^��]�����������U���8�H�A ]�����������������U���8�H�I(]�����������������U���8�H��  ]��������������U���8�H��   ]��������������U���8�H��  ]��������������U���8�H��  ]��������������U���8�H�A$��V�U�WR�Ћ�8�Q�u���BV�Ћ�8�Q$�BDV�Ћ�8�Q$�BLVW�Ћ�8�Q$�JH�E�P�ы�8�B�P�M�Q�҃�_��^��]������U���8�H���  ��V�U�WR�Ћ�8�Q�u���BV�Ћ�8�Q$�BDV�Ћ�8�Q$�BLVW�Ћ�8�Q$�JH�E�P�ы�8�B�P�M�Q�҃�_��^��]���U���8�H���  ]��������������U���<�9��SVW�E�    t�E�P�   ��������/��8�Q�J�E�P�   �ы�8�B$�PD�M�Q�҃��}��8�H�u�QV�ҡ�8�H$�QDV�ҡ�8�H$�QLVW�҃���t)��8�H$�AH�U�R����Ћ�8�Q�J�E�P�у���t&��8�B$�PH�M�Q�ҡ�8�H�A�U�R�Ѓ�_��^[��]���U���8�H�U���  ��VWR�E�P�ы�8�u���B�HV�ы�8�B$�HDV�ы�8�B$�HLVW�ы�8�B$�PH�M�Q�ҡ�8�H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]���������̡�8�H���   ��U���8�H���   V�uV�҃��    ^]�������������U���8�P�]���8�P�B����̡�8�P���   ��U���8�P�R`]�����������������U���8�P�Rd]�����������������U���8�P�Rh]�����������������U���8�P�Rl]�����������������U���8�P�Rp]�����������������U���8�P�Rt]�����������������U���8�P���   ]��������������U���8�P�Rx]�����������������U���8�P���   ]��������������U���8�P�R|]�����������������U���8�P���   ]��������������U���8�P���   ]��������������U���8�P���   ]��������������U���8�P���   ]��������������U���8�P���   ]��������������U���8�P���   ]��������������U���8�P���   ]��������������U���8�P���   ]��������������U���8�P���   ]��������������U���8�P���   ]��������������U���8�P�EPQ��  �у�]� �U���8�P���   ]��������������U���8�P���   ]��������������U���8�P���   ]��������������U��E��t ��8�R P�B$Q�Ѓ���t	�   ]� 3�]� U���8�P �E�RLQ�MPQ�҃�]� U��E��u]� ��8�R P�B(Q�Ѓ��   ]� ������U���8�P�R]�����������������U���8�P�R]�����������������U���8�P�R]�����������������U���8�P�R]�����������������U���8�P�R]�����������������U���8�P�R]�����������������U���8�P�E�R\P�EP��]� ����U���8�E�P�B ���$��]� ���U���8�E�P�B$Q�$��]� �����U���8�E�P�B(���$��]� ���U���8�P�R,]�����������������U���8�P�R0]�����������������U���8�P�R4]�����������������U���8�P�R8]�����������������U���8�P�R<]�����������������U���8�P�R@]�����������������U���8�P�RD]�����������������U���8�P�RH]�����������������U���8�P�RL]�����������������U���8�P�RP]�����������������U���8�P���   ]��������������U���8�P�RT]�����������������U���8�P�EPQ��  �у�]� �U���8�P���   ]��������������U���8�P���   ]��������������U���8�P�RX]����������������̡�8�P���   ��U���8�P���   ]��������������U���8�P���   ]��������������U���8�P���   ]��������������U���8�P���   ]�������������̡�8�P���   ��U���8�P���   ]�������������̡�8�P���   ���8�P���   ���8�P���   ��U���8�H���   ]��������������U���8�H��   ]��������������U���8�H�U�E��VWRP���  �U�R�Ћ�8�Q�u���BV�Ћ�8�Q�BVW�Ћ�8�Q�J�E�P�у�_��^��]������������U���8�H���  ]��������������U���8�P(�BPVW�}�Q�]���E�$�Ѕ�tM��8�G�Q(�]�E�BPQ���$�Ѕ�t,��8�G�Q(�]�E�BPQ���$�Ѕ�t_�   ^]� _3�^]� ����U���8�P(�BTVW�}����$���Ѕ�tE��8�G�Q(�BT�����$�Ѕ�t(��8�G�Q(�BT�����$�Ѕ�t_�   ^]� _3�^]� U��VW�}W��� �����t8�GP���������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U��VW�}W��� �����t8�GP��������t)�O0Q��������t��HW���������t_�   ^]� _3�^]� ������������U���8�} �P(�R8��P��]� ����U���8�P�BdS�]VW��j ���Ћ�8�Q�����   h�+��h�  V�Ћ�8�����Eu�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћ�8�Q(�BHV���Ѕ�t ��8�Q(�E�R VP���҅�t�   �3��EP��j����_��^[]� ����U���V�E���MP�K���P���#�����8�Q�J���E�P�у���^��]� ���h9Ph�����  ���������������U��Vh9h�   h�������  ����t���   ��t�MQ����^]� 3�^]� �U��Vh9h�   h������  ����t���   ��t�MQ����^]� 3�^]� �U��Vh9h�   h�����F�  ����t ���   ��t�M�EQ�����$��^]� 3�^]� ��������U��Vh9h�   h�������  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh9h�   h������  ����t���   ��t�MQ����^]� 3�^]� �U��Vh9h�   h�����f�  ����t ���   ��t�MQ����3҅���^��]� 3�3҅���^��]� ���������������h9h�   h����  ����t���   ��t��3��������U��h9h�   h���ٿ  ����t���   ��t]��]���̋�3ɉH��H�@   �������������U��ыM��tK�E��t��8���   P�B@��]� �E��t��8���   P�BD��]� ��8���   R�PD��]� �����U���8�P@�Rd]�����������������U���8�P@�Rh]�����������������U���8�P@�Rl]�����������������U���8�P@�Rp]�����������������U���8���   ���   ]�����������U���8���   ���   ]����������̡�8�P@�Bt����̡�8�P@�Bx�����U���8�P@�R|]����������������̡�8�P@���   ���8���   �Bt��U���8�P@���   ]�������������̡�8�P@���   ��U���8�P@���   ]��������������U���8�P@���   ]��������������U���8�P@���   ]��������������U���8�P@���   ]��������������U���8V��H@�QV�ҋM����t��#�����8�Q@P�BV�Ѓ�^]� �̡�8�PH���   Q�Ѓ�������������U���8�P@�EPQ�JL�у�]� ���̡�8�P@�BHQ�Ѓ����������������U���8�P@�EP�EP�EPQ�J�у�]� ������������U���8�P@�EPQ�J�у�]� ����U���8�P@�EP�EPQ�J�у�]� U���8�P@�EPQ�J �у�]� ����U���8���   �R]��������������U���8���   �R]��������������U���8���   �R ]��������������U���8���   ���   ]�����������U���8���   ��D  ]�����������U���8�E���   �E ���   P�E���$P�EP�EP�EP��]� ���������U���8���   ���   ]����������̡�8���   �B$���8�H@�Q0�����U���8�H@�A4j�URj �Ѓ�]����U���8�H@�A4j�URh   @�Ѓ�]�U���8�H@�U�E�I4RPj �у�]�̡�8�H|�������U��V�u���t��8�Q|P�B�Ѓ��    ^]��������̡�8�H|�Q �����U��V�u���t��8�Q|P�B(�Ѓ��    ^]��������̡�8�H@�Q0�����U��V�u���t��8�Q@P�B�Ѓ��    ^]���������U���8�H@���   ]��������������U��V�u���t��8�Q@P�B�Ѓ��    ^]��������̡�8�PH���   Q�Ѓ�������������U���8�PH�EPQ��d  �у�]� �U���8�H �IH]�����������������U��}qF uHV�u��t?��8���   �BDW�}W���Ћ�8�Q@�B,W�Ћ�8�Q�M�Rp��VQ����_^]����������̡�8�P@�BT�����U���8�P@�RX]�����������������U���8�P@�R\]����������������̡�8�P@�B`�����U���8�H��T  ]��������������U���8�H@�U�A,SVWR�Ћ�8�Q@�J,���EP�ы�8�Z��h��hE  �΋���2  Ph��hE  ����2  P��T  �Ѓ�_^[]���̡�8�PD�BQ�Ѓ���������������̡�8�PD�BQ�Ѓ���������������̡�8�PD�BQ�Ѓ����������������U���8�PX��Q�
�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ���������U���8�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U���8�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U���8�PX��`VWQ�J�E�P�ы��E���   ���_^��]� �������������U���8�PX�EPQ�J�у�]� ����U���8�PX�EPQ�J�у�]� ����U���8�PX�EPQ�J�у�]� ����U���8�PX�EPQ�J�у�]� ����U���8�PX�EPQ�J$�у�]� ����U���8�PX�EPQ�J �у�]� ����U���8�PD�EP�EPQ�J�у�]� U���8�HD�U�j R�Ѓ�]�������U���8�H@�AV�u�R�Ѓ��    ^]��������������U���8�HD�	]��U���8�H@�AV�u�R�Ѓ��    ^]��������������U���8�HD�U�j R�Ѓ�]�������U���8�H@�AV�u�R�Ѓ��    ^]��������������U���8�U�HD�Rh2  �Ѓ�]����U���8�H@�AV�u�R�Ѓ��    ^]��������������U���8�U�HD�RhO  �Ѓ�]����U���8�H@�AV�u�R�Ѓ��    ^]��������������U���8�U�HD�Rh'  �Ѓ�]����U���8�H@�AV�u�R�Ѓ��    ^]�������������̡�8�HD�j h�  �҃�����������U���8�H@�AV�u�R�Ѓ��    ^]�������������̡�8�HD�j h:  �҃�����������U���8�H@�AV�u�R�Ѓ��    ^]��������������U���3��E��E���8���   �R�E�Pj�����#E���]�̡�8�HD�j h�F �҃�����������U���8�H@�AV�u�R�Ѓ��    ^]�������������̡�8�HD�j h�_ �҃�����������U���8�H@�AV�u�R�Ѓ��    ^]��������������U��E����u��]� �E���8�E�    ���   �R�E�Pj������؋�]� ̡�8�PD�B$Q�Ѓ���������������̡�8�PD�B(Q�Ѓ���������������̡�8�PD�BQ�Ѓ���������������̡�8�PD�B(Q�Ѓ���������������̡�8�PD�BQ�Ѓ���������������̡�8�PD�B(Q�Ѓ���������������̡�8�PD�BQ�Ѓ���������������̡�8�PD�B(Q�Ѓ���������������̡�8�PD�BQ�Ѓ���������������̡�8�PD�B(Q�Ѓ���������������̡�8�PD�BQ�Ѓ���������������̡�8�PD�B(Q�Ѓ���������������̡�8�PD�BQ�Ѓ���������������̡�8�PD�B(Q�Ѓ���������������̡�8�PD�BQ�Ѓ���������������̡�8�PD�B(Q�Ѓ���������������̡�8�PD�BQ�Ѓ���������������̡�8�PD�B(Q�Ѓ���������������̡�8�PD�BQ�Ѓ����������������U���8�E�PH�B���$Q�Ѓ�]� ���������������U���8�PH�EPQ���   �у�]� �U���8�PH�EPQ���  �у�]� �U���8�PH�EPQ���  �у�]� �U���8�PH�EP�EPQ��  �у�]� �������������U���8�PH�EP�EPQ��  �у�]� ������������̡�8�PH���  Q�Ѓ�������������U���8�PH�EPQ���  �у�]� ̡�8�PH���   j Q�Ѓ�����������U���8�PH�EPj Q���   �у�]� ��������������̡�8�PH���   jQ�Ѓ�����������U���8�PH�EPjQ���   �у�]� ��������������̡�8�PH���   jQ�Ѓ����������U���8�PH�EPjQ���   �у�]� ���������������U���8�PH�EP�EPQ���   �у�]� �������������U���8�PH�EP�EPQ���   �у�]� ������������̡�8�PH���   Q�Ѓ�������������U���8�PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP���@���������t�E��8�QH���   PVW�у���_^]� �����U��EVW���MPQ�L���������t�M��8�BH���   QVW�҃���_^]� ̡�8�PH���   Q�Ѓ������������̡�8�PH���   Q�Ѓ�������������U���8�PH�EPQ���   �у�]� �U���8�PH�EPQ���   �у�]� �U���8�PH�EP�EPQ��8  �у�]� �������������U���8�PH�EP�EPQ��   �у�]� ������������̡�8�PH���  Q�Ѓ������������̡�8�PH���  Q�Ѓ������������̡�8�PH���  Q�Ѓ������������̡�8�PH��  Q�Ѓ������������̡�8�PH��  Q�Ѓ�������������U���8�PH�EP�EPQ��  �у�]� �������������U���8�PH�EP�EP�EPQ��   �у�]� ���������U���8�PH�EP�EP�EP�EPQ��|  �у�]� �����U���8�PH�EPQ��  �у�]� ̡�8�PH��T  Q�Ѓ�������������U���8�PH�EP�EPQ��  �у�]� �������������U���8�PH�EPQ��8  �у�]� �U���8�PH�EPQ��<  �у�]� �U���8�PH�EPQ��@  �у�]� �U���8�PH�EP�EP�EPQ��D  �у�]� ��������̡�8�PH��L  Q��Y��������������U���8�PH�EPQ��H  �у�]� ̡�8V��H@�Q,WV�ҋ�8�Q��j �ȋ��   h�  �Ћ�8�QH�����   h�  V�Ѓ���
��t_3�^Ë�_^�̡�8�P@�B,Q�Ћ�8�Q��j �ȋ��   h�  �������U���8�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U���8�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U���8�PH�EP�EP�EPQ��   �у�]� ��������̡�8�HH��  ��U���8�HH��  ]��������������U���8�E�PH��$  ���$Q�Ѓ�]� �����������̡�8�PH��(  Q�Ѓ�������������U���8�PH�EP�EPQ��,  �у�]� �������������U���8�E�PH�EP�E���$PQ��0  �у�]� ���̡�8�PH���  Q�Ѓ������������̡�8�PH��4  Q�Ѓ������������̋��     �������̡�8�PH���|  jP�у���������U���8�UV��HH��x  R��3Ƀ������^��]� ��̡�8�PH���|  j P�у��������̡�8�PH��P  Q�Ѓ������������̡�8�PH��T  Q�Ѓ������������̡�8�PH��X  Q�Ѓ�������������U���8�PH��Q��\  �E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����̡�8�PH��`  Q�Ѓ�������������U���8�PH�EPQ��d  �у�]� �U���8�E�PH��h  ���$Q�Ѓ�]� ������������U���8�E�PH��t  ���$Q�Ѓ�]� ������������U���8�E�PH��l  ���$Q�Ѓ�]� ������������U���8�PH�EPQ��p  �у�]� �U���8�PH�EP�EP�EP�EPQ���  �у�]� �����U���8�PH�EP�EP�EP�EP�EP�EPQ���  �у�]� �������������U���8�E�HH�U �ER�UP�E���$R�UP���   R�Ѓ�]������������U��U�E��8�HH�E���   R�U���$P�ERP�у�]����������������U���E�M��'��� �M;�|�M;�~��]�����������U���8�PH�E���   Q�MPQ�҃�]� ������������̡�8�PH���   Q��Y�������������̡�8�PH���   Q�Ѓ������������̡�8�PH���   Q��Y��������������U���8�PH�EP�EPQ���   �у�]� �������������U���8�PH�EP�EP�EP�EP�EPQ���  �у�]� ̡�8�PH��t  Q��Y�������������̋�� �+�@    ���+��8�Pl�A�JP��Y��������U���8V��Hl�V�AR�ЋE����u
�   ^]� ��8�Ql�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uË�8�QlP�B�Ѓ�������U���8�Pl�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U��U�E��8�HH�ER�U���$P���  R�Ѓ�]����U���8�HH���  ]��������������U���8�HH���  ]��������������U��U0�E(��8�HH�E$R�U ���$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�,]������������U���8�HH���  ]��������������U���8�E�PH�EP���$Q���  �у�]� ��������U���SV����  �؅ۉ]���   �} ��   ��8�HH��p  j h�  V�҃����E�u
^��[��]� �MW3��}���  ����   �]��I �E�P�M�Q�MW�_�  ��tc�u�;u�[�I ������u�E�������L�;Ht-��8�Bl�S�@����QR�ЋD������t	�M�P�C�  ��;u�~��}��M���}��
�  ;��r����]�_^��[��]� ^3�[��]� ����������U�����8SV�ًHH��p  j h�  S�]��ҋ�����u
^3�[��]� �E��u��8�HH���  �'��u��8�HH���  ���uš�8�HH���  S�ҋȃ��ɉEt�W���  ��8�HH���   h�  S3��҃����  ���_�u����    ��8�Hl�U�B�IWP�ы�������   ��8�F�J\�UP�A,R�Ѓ���t�K�Q�M���  ��8�F�J\�UP�A,R�Ѓ���t�K�Q�M���  �E��;Pt&�F��8�Q\�J,P�EP�у���t	�MS��  ��8�v�B\�M�P,VQ�҃���t�M�CP�s�  ��8�QH�E����   �E�h�  P�����у�;�����_^�   [��]� ������U���8�HH���   ]�������������̡�8�PH���   Q��Y��������������U���8�HH���  ]��������������U���8��P���   V�uW�}���$V�����E������At���E������z����؋�8�Q�B,���$V����_^]����������������U���0���8�U�V�u�U��]�W�P�}���   �E�PV�M�Q����� �@�@�E�����E��Au�����������z���������������z�����������Au������������z)���١�8�]��ɋ��]��]��P�RH�E�PV��_^��]���������Au������������������U���8�HH�]��U���8�H@�AV�u�R�Ѓ��    ^]�������������̡�8�HH�h�  �҃�������������U���8�H@�AV�u�R�Ѓ��    ^]��������������U���8�HH�Vh  �ҋ�������   �EPh�  ��������t]��8�QHj P���   V�ЋMQh(  �V�������t3��8�JH���   j PV�ҡ�8���   �B��j j���Ћ�^]á�8�H@�QV�҃�3�^]�������U���8�H@�AV�u�R�Ѓ��    ^]��������������U���8�HH�Vh�  �ҋ�����u^]á�8�HH�U�E��  RPV�у���u��8�B@�HV�у�3���^]�������U���8�H@�AV�u�R�Ѓ��    ^]��������������U���8�HH�I]�����������������U���8�H@�AV�u�R�Ѓ��    ^]��������������U���8�PH�EPQ���  �у�]� �U���8�PH�EPQ���  �у�]� ̡�8�PH���  Q�Ѓ�������������U���8�HH���  ]��������������U���8�E�HH�U0�E,R�U(P�E$R�U P�ER�U���\$�E�$P��P  R�Ѓ�,]������������̡�8�PH���  Q�Ѓ�������������U���8�PH�EP�EPQ���  �у�]� ������������̡�8�PH��  Q�Ѓ�������������U���8�PH�EP�EP�EPQ���  �у�]� ��������̡�8�PH���  Q�Ѓ������������̡�8�PH���  Q�Ѓ�������������U���8�PH�EPQ��  �у�]� �U���8�PH�EPQ��  �у�]� ̋������������������������������̡�8�HH���  ��U���8�HH���  ]��������������U���8�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ���������U���8�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ��������̡�8�PH��,  Q�Ѓ�������������U���8�PH�EPQ��X  �у�]� ̡�8�PH��\  Q�Ѓ�������������U���8�HH��0  ]��������������U���8��W���HH���   j h�  W�҃��} u�   _��]� Vh�  �������������   ��8�HH���   j VW�҃��M��  ��8�P�E�R0Ph�  �M����E��8�P�B,���$h�  �M��Ћ�8�Q@�J(j �E�PV�у��M��  ^�   _��]� ^3�_��]� �����U��S�]�; VW��u7��8�U�HH���   RW�Ѓ���u��8�QH���   jW�Ѓ���t�   �����   ��8�QH���   W�Ѓ��} u(��8�E�QH�M���  P�ESQ�MPQW�҃��B�u��t;��8�U�HH�ER�USP���  VRW�Ћ�8���   �B(�����Ћ���uŃ; u��8�QH���   W�Ѓ���t3���   ���Wu1��8�QH���   �Ћ�8�E�QH���   PW�у�_^[]� ��8�BH���   �у��} u0��8�M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� ��8�QH�h  �Ћ؃���u_^[]� ��8���   �u�Bx���Ћ�8���   P�B|���Ѕ�tU��8�E�QH�MP�Ej Q���  VPW�у���t��8���   �ȋBHS�Ћ�8���   �B(���Ћ���u�_^��[]� ��������������U��E��V��u��8�HH���  �'��u��8�HH���  ���u��8�HH���  V�҃���u3�^]� P�EP���>���^]� ���������U���D��8�HH���   S�]VWh�  S�ҋ��8�HH���   3�Wh�  S�u܉}��҃�;��E�}�}��}��p
  ��8���   �B����=�  ��8�  �QH���   Wh:  S�Ћ�8�QH�E����   h�  S�Ћ�8�QHW�����   h�  S�uԉ}��Ћ�8�QH�E苂  S�Ћ�8�QH�EЋ��  S�Ѓ�(���E��E��+�}   �M���M�MЅ�tMj�W�0�  ���t@�@�Ẽ|� �4�~����%�������;�u/���O�  ;E�~�E؋���  E���E�;Pu�E���E��E���;}�|��}� tv�u�j S�����������  ���������tV�������}�;�uK��8�H���  �4�h�+��h�  V�҃����E��k  �M�PVP����P��  ����}ܡ�8�H���  �4�h�+��h�  V�҃����E��   �M�3�;�t;�tVQP��} ���E�;�~-��8�Qh�+��h�  P���   �Ѓ�;ǉE���  ��8�E��QH��  j�PS�у�����  �u�;�tjS�����������  ��������E���}��8�BH���   Wh�  S�у�3�9}ԉE�}���  �}���}ȋMЅ��p  �U�j�R�8�  ����\  �M̍@�|� ���]�~����%�������9E��  ����  �E�3�3�9C�E܉M���   ��I �����������t{�]��}������������ϋ9�<��}����҉��y�]��|��]������z�<��y�]��|��]������z�<��I�}��]������M��}ȃ��������M؃�;K�M��b������E��O  �+U�j��PR�M��c�  �M�v���E�3�+��U��E����	��$    ���E�;E���   �}� �U����E�t6�U�@�U�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�M��E�;]؍@�E��Ћ��P�Q�P�Q�P�Q�P�Q�@�A}c�UȋE�9�uX�ȋL�����������w4�$�H�U����4�"�M����t��U����t�
�M����t�M���;]�|��E�����;]؉M������U�;U��  �U�R�Q5���E�P�H5���M�Q�?5����_^3�[��]Ë�M�3�;G�Å���   �E�v�ЋW��R�ы��Q�P�Q�P�Q�P�Q�P�I�H�O��I�M�ы�P�Q�P�Q���ۉP�Q�P�Q�P�I�H��@�E�ЋU�Lv�ʋ��P�Q�P�Q�P�Q�P�Q�@�At8�G�U�@�ʋU�Lv	�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��w��U��@�ʋU���v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��w��U����@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�7����t?�G�U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�w�����O�E�����;EԉE��}�������U�R�'3���E�P�3�����$  ���   �B����=  �  ��8�QH���   j h(  S�Ћ�8�QH�����   h(  S�ЋЃ�3��҉U�~#���ǅ�t�|� t�4N��tN���;�|�u��u܋�8�Q���  �4v�h�+��hK  V�Ѓ����E���   �M��t��tVQP��w ���u؋�8�Q���  �h�+��hP  V�Ѓ����E�tP��t��tVWP�w ���M����+�8�RH��PQ�E���   S�Ѓ���u�M�Q��1���U�R��1����_^3�[��]á�8�HH���   j h�  S�҉E���8�HH���   j h(  S��3�3���3�9]؉E��}ĉ]��N  �U���    �څ��+  ���E�    ��   �U�<��v��   ����U��:��\:�Y�\:�Y�\:׉Y�Z�Y�R�Q�U��\�E��Y�\�T���Y�Z�Y�Z�Y�Z�Y�R�]��Q�U�����������;�|��}ă|� �w   �U��Eԍ8�I�ʋU�v���A�B�A�B�A�B�A�B�I�J�E���ЋE���v�Ћ��A�B�A�B�A�B�A�B�I�J�U���<ډ}ă�;]؉]�������M�3�3�;�~"�U����$    �d$ �t���   ��;�|�U�R��/�����E�P��/����_^�   [��]Ë�lw����������U��U��t�M��t�E��tPRQ�0u ��]������������U��E� �M+]� ���������������U��V��V��+��8�Hl�AR�Ѓ��Et	V�2������^]� ���������̡�8�P�BVj j����Ћ�^���������U���8�P�E�RVj P���ҋ�^]� U���8�P�E�RVPj����ҋ�^]� ��8�P�B�����U���8�P���   Vj ��Mj V�Ћ�^]� �����������U���8�P�EPQ�J�у�]� ����U���8�P�EPQ�J�у������]� �������������U���8�P�E�RtP�ҋ�8���   P�BX�Ѓ�]� ���U���8�P�E�Rlh#  P�EP��]� ���������������U���8�P�E�RlhF  P�EP��]� ���������������U���8�P�E�RtP�ҋ�8���   �M�R`QP�҃�]� ���������������U���8�P���   ]��������������U���8�P�E���   P�҅�u]� ��8���   P�B�Ѓ�]� ��������3��������������̃��� ���������̸   � ��������3�� ����������̸   � ��������3�� ����������̸ }  � �������̃��� ���������̃��� ���������̃��� ����������U��E�     ]� ���� ����������U����   V�u��u3�^��]�h�   ��@���j P�m �M�Eh�   ��@���R��@����MPQjǅD���PJ��`����E��N�E�`%�E� �E��u�E� O�E��u�8���� ^��]����������������U����   V�u��u3�^��]�h�   ��@���j P�m �M�Uh�   ��@���P��@����M�U��UQRjǅD���PJ��`����E��N�E� �E�`%�E� O�E��u�E�O�E��u�E��u�S7���� ^��]������������U���8�P�B<��   V�uW���Ѕ��}tj VW�C������u_^��]�h   ������j Q�3l �U�E�MRj j PQ������R��O���Mh   ������PQWj�E���E��6����8_^��]���������U���8�P�B<��   V�uW���Ѕ��}tj VW�������u_^��]�h   ������j Q�k �U �E�MRj j PQ������R�7O���U�Eh   ������QRWj�E��E���6����8_^��]���������̋�`�����������U���8�PT�EP�EPQ�J�у�]� U���8�PT�EPQ�J�у�]� ����U���8�PT�EPQ�J�у�]� ����U���8�PT�E�R<��PQ�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U���8�HT�]��U���8�H@�AV�u�R�Ѓ��    ^]�������������̡�8�HT�hG  �҃�������������U���8�H@�AV�u�R�Ѓ��    ^]��������������U���V�u�W�}�����Dz�F�_����D{:�F����$�J� �G��$�]��:� �E���������D{_�   ^��]�_3�^��]���������U���VW�M�������E���}t-��8�Q4P�B�Ѓ����M�u�����_3�^��]Ë�R(���8�H0�QW�҃����M�tԋ�R Q�MQ���ҋ��8�P�B �M��Ѓ��t��8�Q0�Jx�E�PW�у��M�����_��^��]�������U���8�P�B VW�}�����=NIVb��   ��   =TCAbtR=$'  t6=MicM��   ��8�Q���   j hIicM���ЋWP�B����_^]� ��BW����_�   ^]� ��8�Q���   j hdiem���ЋWP�B����_^]� =INIb��   �~ u���B���F   ��_^]� �~ t���B����_^]� =atniDt5=ckhct=ytsdu?��B����_�F    3�^]� ��B����_^]� �A3��_3�^]� =cnys����_3�^]� ������V���4,��8�H0�Vh '�҉F���F    ��^�����V��F���4,t��8�Q0P�B�Ѓ��F    ^�����̡�8�P0�A���   P�у����������U���8�P0�E�I���   PQ�҃�]� �������������̡�8�I�P0���   Q�Ѓ���������̡�8�P0�A���   j j j j j j j j j4P�у�(������̡�8�P0�A���   j j j j j j j j j;P�у�(�������U���8�P0�E�IPQ���   �у�]� ��������������U����E V��P�M�������8�E�Q�R4Ph8kds�M��ҡ�8�E     �H0���   �U R�U�E�P�Ej R�UP�ER�UP�FRj2P�ыu ��(�M��X�����^��]� ��������������̡�8�I�P0���   Q�Ѓ����������U��V��F��u^]� ��8�Q0�M ���   j j j j j Q�Mj QjP�ҡ�8�H0�U�E���   R�UP�ER�UP�Fj RP�у�D^]� ���̋A��uË�8�Q0P�B�Ѓ������̋A��u� ��8�Q0P�B�Ѓ�� �U��Q����u�E�    �P��]� �E�H� V�5�8�v0Q�MQP���   R�U�R�Ћu�    �F    ��8���   j P�BV�Ћ�8���   �
�E�P�у�$��^��]� �������U���8�P0�E�I�RPQ�҃�]� �U��A��t)��8�Q0�M���   j j j j j j Qj jP�҃�(]� ���������U��Q��u3�]� �E�H� V�5�8�v0Q�MQPR�V�҃�^]� ����������U��Q��u3�]� �E�H� V�5�8�v0QP���   R�Ѓ�^]� �����������U��Q��u3�]� �E�H� V�5�8�v0Q�MQPR�V\�҃�^]� ����������U��y u3�]� V�u�W�}�؉��ډ��8�P4�A�JhWVP�ы�ډ����ى_^]� �����U��A��u]� ��8�Q4�M�RhQ�MQP�҃�]� ����U��A��u]� ��8�Q4�M�RpQ�MQP�҃�]� ����U��y u3�]� V�u�W�}�؉��ډ��8�P4�A�JpWVP�ы�ډ����ى_^]� �����U���$VW��htniv�M��i�����8�P�E�R4Phulav�M��ҡ�8�P�B4hgnlfhtmrf�M��Ћ�8�E�Q�R4Phinim�M��ҡ�8�P�E�R4Phixam�M��ҡ�8�P�E�R4Phpets�M��ҡ�8�P�E�R4Phsirt�M��ҋE =  ��}$u�����t.��8�QP�B4h2nim�M��Ћ�8�Q�B4Wh2xam�M��ЋU�M�QR�E�P���K�����8���   P�B8�Ћ�8���   �
���E�P�у��M�����_��^��]�  ��������������U���$V��htlfv�M������E��8�P�B,���$hulav�M��Ћ�8�E,�Q�R4Phtmrf�M����E��8�P�B,���$hinim�M����E��8�Q�B,���$hixam�M����E$��8�Q�B,���$hpets�M��Ћ�8�ED�Q�R4Phsirt�M��������E0��������Dzw���]8����Dzm�؋�8�E@�Q�R4Phdauq�M��ҋM�E�PQ�U�R���������8���   P�B8�Ћ�8���   �
���E�P�у��M��,�����^��]�@ �١�8�P�B,���$h2nim�M����E8��8�Q�B,���$h2xam�M����V�����U���$V��hgnrs�M������E��8�E��E�   �Q���   �E�Pj�M��ҡ�8���   ��U�R�ЋM��8�M����E�   �B���   �M�Qj�M��ҡ�8���   ��U�R�ЋU���M�QR�E�P���������8���   P�B8�Ћ�8���   �
���E�P�у��M��
�����^��]� �U���$V��hCITb�M�������8�P�E�R8PhCITb�M��ҡ�8�P�E�R4Phsirt�M��ҡ�8�P�E�R4Phulav�M��ҋM�E�PQ�U�R��������8���   P�B8�Ћ�8���   �
���E�P�у��M��Y�����^��]� U��E��Vj ��P�M�Q�M赑���UPR���)������8�H�A�U�R�Ѓ���^��]� ����������U��E,��UPj ���T$�$htemf�E$�� �\$�E�\$�E�\$�E�$R�O���]�( �����������U��E,��Pj ���T$�U�$hrgdf�E$�� ��$����$�����\$�E�����\$�M���\$�E�$R�����]�( ���U��E,��Pj ���T$�U�$htcpf�E$�� ��'�����\$�E���\$�}�\$�E�$R����]�( ���������������U��Q��u3�]� �E�E�H� V�5�8�v0Q�M Q�M���\$�E�$QPR�V(�҃�$^]� ������U��Q��u3�]� �E�H� V�5�8�v0Q�MQPR�V,�ҋU3Ƀ�9M^���
]� �������������U��Q��u3�]� �E�H� V�5�8�v0Q�MQPR�V,�҃�^]� ����������U��Q��u3�]� �E�H� V�5�8�v0Q�MQPR�V0�҃�^]� ����������U��SVW���W��t$�E�H�5�8�^0� �uQVP�C0R�Ѓ���u	_^3�[]� �W��t��E�H� ��8�[0Q�NQPR�S0�҃���t̋W��tŋE�H� �=�8�0Q��VP�G0R�Ѓ���t�_^�   []� ��U��Q��u3�]� �E�H� V�5�8�v0Q�MQ�MQPR�V<�҃�^]� ������U��QV3���Wu3��,�E�H� �5�8�v0Q�MQPR�V,��3Ƀ�9M�������8�M�B�P0VQ�M�ҋ�_^]� ����U��A��Vu3��"�M�Q�	�5�8�v0R�URQP�F,�Ѓ�����8�Q�E�M�R4PQ�M�ҋ�^]� ���������������U��A����Vu3��"�M�Q�	�5�8�v0R�U�RQP�F0�Ѓ�����8�E��Q�E�M�R,���$P�ҋ�^��]� �����U�����V���U��V�U����]�Wt$�E�H� �=�8�0Q�M�QPR�W0�҃���u
_3�^��]� �V��t�E�H� �=�8�0Q�M�QPR�W0�҃���tˋV��tċE�H� �5�8�v0Q�M�QPR�V0�҃���t���8�P�M�RH�E�PQ�M��_�   ^��]� �����������U��� ��A���U�V�U��]�Wu3��&�M�Q�	�5�8�v0R�U�R�U�RQP�F<�Ѓ����E����}t��8�Q�RH�M�QP���ҋE���t��8�E��Q���$P�B,����_��^��]� U���8�P�E���   Vj ��MP�ҋM$�U Q�MR�Uj Q�MR�UQPR���o���^]�  ����������U���8��P�E���   V���$��MP���E8�E@�M,�Uj P���\$�E0�$Q�E$�� �\$���E�\$�E�\$�$R�K���^]�< ������U���8��P�E���   V���$��MP����Ej j ���T$���$htemf�E$�� �\$�E�\$�E�\$�$P�����^]�$ �����������U���8��P�E���   V���$��MP���E$�Ej �� �\$���E�\$�E�\$�$P�C���^]�$ ��������������U���8��P�E���   V���$��MP����j j ���T$�E�$htcpf�E$�� ��'�������\$�E���\$�}�\$�$P����^]�$ ���������������U���8�� V��H�A�U�R�ЋM�E��Qj �U�RP�M�Q�M������UPR���������8�H�A�U�R�Ћ�8�Q�J�E�P�у���^��]� ������������U���dV��M�蟇����8�Q���   P�EP�M�Q�M��P�M��)����M��a���j j �E�P�M������MPQ��������8���B�P�M�Q�҃��M��&����M�������^��]� �����U���P��E����]���VW�}��t��8�Q���$P���   �����]����8�U��UЍE��]ȋQ�M���   PQ�E�P���ҋ�M��P�U�H�M�P�U�H�M��P�F���U�u_^��]� �M�E�Q�	�5�8�v0R�U R���\$�U��E��$RQP�F(�Ѓ�$_^��]� ���������������U���0�E���M�u��8�H���   �҅�u��]� SVW���o����htlfv�MЉu������E�}��8�X�U�����$��i �]��G�$��i �}�S,�M��$hulav�ҡ�8�P�B4hmrffhtmrf�M��Ћ}���8�M�Y���$�i �]��G�$�i �}�S,�M��$hinim�ҋ}���8�M�X���$�Yi �]��G�$�Ki �}�S,�M��$hixam�����8�P�B,���$hpets�M��Ћ�8�Q�B4j hdauq�M��Ћ�8�Q�B4Vhspff�M��Ћ�8�E �Q�R4Phsirt�M��ҋM�E�PQ�M��U�R�n�����8���   P�B8�Ћ�8���   �
���E�P�у��M�����_��^[��]� U��E����V��u��8�H���   �҅�u^��]� ����m���E�F��u3��"�M�Q�	�5�8�v0R�U�RQP�F0�Ѓ����E����'�M������\$�M��$��  ��M��P�Q�P�Q�@�A��^��]� ����������U���0���8�]�V���M�]�P���   �E�PQ�M�E�P�ҋ�P�M��Hj �U�P�E P�M��MQ�M�U��UR�U�E�PQR������^��]� ���������������U�����UV�]���E�P�]��ERP������8�Q�M�R@���E�PQ�M�ҋ�^��]� ����������U��A��u]� �M�Q�	V�5�8�v0Rj j j j j j Qj1P���   �Ѓ�(^]� ���������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��A��u]� ��8�Q0�M���   j j j j j j j Qj-P�҃�(]� �����U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj j j Q�MQj j j)P�ҋE���(��]� ��U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj j Q�Mj Qj j j)P�ҋE���(��]� ��U��A��u]� ��8�Q0�M���   j j j Q�MQ�MQ�Mj Qj/P�҃�(]� ���������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj'P�ҋE���(��]� ������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj,P�ҋE���(��]� ������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�MQ�MQjP�ҋE���(��]� ����������U���8�P0�E�I���   j j j P�EP�EP�Ej Pj.Q�҃�(]� ��������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj:P�ҋE���(��]� ������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj*P�ҋE���(��]� ������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj	P�ҋE���(��]� ��������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj
P�ҋE���(��]� ��������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��A��u]� ��8�Q0�M���   j j j Q�MQ�MQ�Mj QjP�҃�(]� ���������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj>P�ҋE���(��]� ������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� �M�Q�	V�5�8�v0R�Uj j j j R�URQjP���   �Ѓ�(^]� �����������U����ESVW�M�P�M��I  �MQ�U�R�M��XI  ��tm�}��E��tN��8���   P�BH�ЋM��I����tQ�W�7��8�[0R�U�j j j j RP���   VjQ�Ѓ�(��t"�MQ�U�R�M���H  ��u�_^�   [��]� _^3�[��]� ��������������U��A��u]� �M�Q�	V�5�8�v0Rj j j j j j QjP���   �Ѓ�(^]� ���������������U��Q�A��u��]� ��8�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� ��8�Q0�M�RDQ�MQ�MQP�҃�]� U��A��u]� ��8�Q0�M�RHQ�MQ�MQ�MQ�MQ�MQP�҃�]� ���̋A��uË�8�Q0P�BX�Ѓ�������U��A��u]� ��8�Q0�M�RLQ�MQP�҃�]� ����U��A��u]� ��8�Q0�M�RP��   �QP�҃�]� ��U��A��u]� ��8�Q0�M�RPQP�҃�]� ��������U��A��u]� ��8�Q0�M�RTQ�MQ�MQ�MQP�҃�]� ������������U���8V�u�VW���H4�R�ЋE�F    �~�H� ��8�R0Q�MQ���   VP�GP�у�3҅��F_^��]� ���U��A��u]� ��8�Q0�M���   j j j j j Qj j jP�҃�(]� �����U��E��u]� �@    �@�I��8�R0P�EPQ���   �у�]� ������̡�8�I�P0���   j j j j j j j j j0Q�Ѓ�(�������U��E��u��8� ��8�R0�I�R@V�uVP�EPQ�҃�^]� �����������U���8�P0�E�I�RdP�EP�EP�EP�EPQ�҃�]� �U���8�P0�E�I�RpP�EP�EP�EP�EPQ�҃�]� �U��E�P� V�5�8�v0R�UR�UR�UR�URP�A�NhP�у�^]� ��������U��E� ��8�R0j j j j j j j P�A���   jP�у�(]� �����������U��E� ��8�R0j j j j j jj P�A���   jP�у�(]� �����������U��E� ��8�R0j j j j j j j P�A���   jP�у�(]� �����������U���V��M������E�H� ��8�R0Q�M�Q���   j j j j j P�Fj8P�ы���(��t�M�U�R�;����M��#�����^��]� ����������U��E�P� V�5�8�v0R�URj j j j j P�A���   j9P�у�(^]� �����U��E�P� V�5�8�v0Rj j j j j j P�A���   j"P�у�(^]� �������U��E�P� V�5�8�v0Rj j j j j j P�A���   j5P�у�(^]� �������U��E�P� V�5�8�v0R�Uj j j j Rj P�A���   j<P�у�(^]� �����U���8�P0�E�I���   j j P�EP�EP�EP�Ej Pj3Q�҃�(]� ������U���8�UVj j j j j R��H0�E�Vj P���   jR�Ћ�8�Q0�E�N�RtPQ�҃�0^]� ��U���8�P0�E�I���   j j j j j j Pj jQ�҃�(]� �������������̡�8�P0�A���   j j j j j j j j jP�у�(�������U���8�P0�E�I���   j j j j j j j PjQ�҃�(]� �������������̡�8�P0�A���   j j j j j j j j j(P�у�(�������U���8�P0�E�I���   j j j j j j P�EPj&Q�҃�(]� ������������U���8�P0�E�I���   j j j j P�EP�Ej Pj+Q�҃�(]� ���������̡�8�P0�A���   j j j j j j j j jP�у�(������̡�8�P0�A���   j j j j j j j j j#P�у�(�������U��QS�]VW�}���M�t��8�P���   j j���Љ�u��t��8�Q���   j j���Љ��8�Q0�E��H�R`VWQ�҃�_^[��]� �U���8�P0�E�I���   P�EP�EPQ�҃�]� �����̡�8�P0�A���   j j j j j j j j j P�у�(������̸   ����������̸   ��������������������������̸   � ��������3�� �����������3���������������� �������������V���4,��8�H0�Vh '�҉F3��F�F���\,�F   ��^�������V��F���4,t��8�Q0P�B�Ѓ��F    ^������U��E�UVj ��MP�EQ3�9MR��Pj �F    ��
Q��������t�~ t
�   ^]� 3�^]� �U��E�A�I��u3�]� ��8�B0Q�H�у�]� ����U���8�P�B S�]V�����=ckhc��   ��   =cksate=TCAb��   ��8�Q���   Wj hdiem���Ћ���BSW���F   �Ѓ~ ��t��t��u3Ƀ���Q���C���_^��[]� �~ tK��B����^[]� �~ t6��������t+�F    ^�   []� =atnit�MQS���/���^[]� ^3�[]� �U��V��~ ��   W�}����   �$��V�E;E��   �r�M;M��   �d�U;U��   �V�E;E��   �H�E;E~@;E��   �5�E;E|-;E~v�&�E;E|;E|g��E;E~;E~X��M;MuN��8�M�B0�V���   j j j j j j j QjR���E��(j���\$�E�$W������F    _^]� �U�U�U�UVV.V=VLV����U��V��~ �  �E W�}�E����   �$� X���]������   �   ���]����A��   �   ���]����A��   �r���]������   �`�E������A��uN��������   �C�E��������u1������A{{�*�E���������E������A�����]����DzU����ء�8�U�H0�F���   j j j j j j j RjP���E �U(��(R���\$�E�$W�S�����F    _^]�$ �I �VW$W6WHWeW~W�W�W������������U���E �E�Uj���\$�E�\$�E�$PR�w���]�  ���U���E �E�Uj���\$�E�\$�E�$PR�G���]�  ���U���E �E�Uj���\$�E�\$�E�$PR����]�  ��̋�3�� �,�H�H�H�������������VW��3�9~��,u��8�H4�V�R�Ѓ��~�~_^����U���8�P4�E�I�RtPQ�҃�]� �U��U��t3�A��8�I0R���   P�ҋ�8�Q0�M���   QP�҃�]� ��8�P0�E�I�R|PQ�҃�]� ������̡�8�P4�A�JP�у������������̡�8�P4�A�JP�у������������̡�8�P4�A�JP�у������������̡�8�P4�A�J|P�у������������̡�8�P4�A���   P�у����������U���8�P4�E�I�RP�EP�EP�EPQ�҃�]� �����U���8�P4�E�I�RP�EP�EP�EPQ�҃�]� �����U���8�P4�E�I�R PQ�҃�]� �U���8�P4�E�I�R$PQ�҃�]� �U���8�P0�E�I���   P�EP�EP�EPQ�҃�]� ��U���8�P4�E�I���   PQ�҃�]� ��������������U���8�P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U���8�P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U���8�P4�E�I�R(PQ�҃�]� �U���8�P4�E�I�R,P�EP�EPQ�҃�]� ���������U���8�P4�E�I�R0P�EPQ�҃�]� ������������̡�8�P4�A�J4P��Y��������������U����UV��EP�M�Q�NR�E�    �E�    ������8�H4�V�AR�Ћ�8�Q0�Rhj �M�Q�M�Q�M�Q�M�QP�F�HQ�҃� �} ^t(�} t(�E��M�;�~<�U��;�}3�E�M�;�~)�U���} u�E��M�;�~�U��;�}�   ��]� 3���]� ��������������U���8�P4�E�I�R8PQ�҃�]� �U���8�P4�E�I�R<PQ�҃�]� �U���8�P4�E�I���   P�EPQ�҃�]� ���������̡�8�P4�A�J@P�у�������������U���8�P4�E�I�RDP�EPQ�҃�]� �������������U���8�P4�E�I�RHP�EPQ�҃�]� �������������U���8�P4�E�I�RLP�EPQ�҃�]� �������������U���8�P4�E�I�RPP�EPQ�҃�]� �������������U���8SV�uW�����   �QV�҃�����   ��8���   �]�QS�҃���SuA��8���   �Q@�ҋء�8���   �Q@V�ҋ�8�Q4�JPSP�GP�у�_^[]� ��8���   �H�у���uD��8���   �H8S�ы�8�؋��   �H@V�ы�8�J4�WSP�AHR�Ѓ�_^[]� h�,h}  ��   ��8���   �BV�Ѓ�����   ��8���   �]�BS�Ѓ���SuC��8���   �B@�Ћ�8���   �؋B8V�Ћ�8�Q4�JLSP�GP�у�_^[]� ��8���   �H�у���uD��8���   �H8S�ы�8�؋��   �H8V�ы�8�J4�WSP�ADR�Ѓ�_^[]� h�,h�  �
h�,h�  ��8�Q��0  �Ѓ�_^[]� �U���8�P4�E�I��  P�EP�EP�EPQ�҃�]� ��U���8�P4�E,P�E(P�E$P�E �IP�E�RTP�EP�EP�EP�EP�EPQ�҃�,]�( �������������U���8�P4�E�I�RXP�EP�EP�EPQ�҃�]� ����̡�8�P4�A�J`P��Y�������������̡�8�P4�A�JdP�у�������������U���8�P4�E�I��   P�EP�EP�EPQ�҃�]� ��U���8�P4�E�I�R\P�EP�EP�EP�EP�EPQ�҃�]� �������������U���8�P4�E�I�RhP�EPQ�҃�]� �������������U��V�u��Wt��؉�}��t��ډ��8�P4�A�JhWVP�у���t��ډ��t��ى_^]� �U��V�u��Wt��؉�}��t��ډ��8�P4�A�JpWVP�у���t��ډ��t��ى_^]� �U���8�P4�E�I�RpP�EPQ�҃�]� �������������U���,V��~ ��   ��8�V�H4�AR�Ѓ} t ��8�Q0�RlP�F�HQ�҃�^��]� ��hARDb�MԉE��E�    �ܼ��P�M�Q�N�U�R������8���   ��U�R�Ѓ��M�����^��]� ������U���8�P4�E�I�RlPQ�҃��   ]� ������������U���8�E�P4�E�I���   P�E���\$�E�$PQ�҃�]� ����������U���8�P4�E�I���   P�EP�EPQ�҃�]� �����̡�8�P4�A���   P�у���������̸   ����������̸   �����������U���8V��H4�V�A$h�  R�Ћ�8�Q4�E�MP�EQ�MP�FQ�JP�у�2�^]� ��������U��U��@R�UR�UR�UR��]� �̸   � ��������3�� ������������ �������������3�� ������������ �������������U���8�P4�E�I�RxP�EP�EP�EPQ�҃�]� �����U���8�P0�E�I�I���   P�EP�EPQ�҃�]� ���U��QS�]VW�}���M�t��8�P���   j j���Љ�u��t��8�Q���   j j���Љ��8�Q4�E��H�RpVWQ�҃�_^[��]� �U��Q��8�P�B SVW�}���3���=INIb�/  �  =SACbvt+=$'  t
=MicM�  ��B$W����_�   ^��[��]� ��R3��E��E�EP�M�Q���҅�t��8�U�H4�E�R�VP�AR�Ѓ�_�   ^��[��]� =ARDb�  ��8�Q���   j j���Ћ�8�Qj �؋��   j���Ћ�8�Qj �E����   j���Ћ�8�Qj �E���   j���ЋM���RWP�EPQS����_�   ^��[��]� ��P����_�   ^��[��]� =NIVbetJ=NPIbt0=ISIbu\�>���Y���P���1���P�G����_�   ^��[��]� ��BW����_^[��]� ��B����_�   ^��[��]� =cnyst_^��[��]� ��8�Q���   j hIicM���ЋWP�B ����_^[��]� �������������U���8�P4�E�I�RTh����h����h����P�EP�Eh����h����h����h����PQ�҃�,]� ������U���V��hYALf�M�躷����8�Q4�JlP�FP�у��M��ܷ��^��]��������V���4,��8�H0�Vh '�҉F���F    ��,�F   ��^��������V��F���4,t��8�Q0P�B�Ѓ��F    ^������U���8�P�B VW�}�����=cksat`=ckhct�MQW��譾��_^]� �Nj j j j j j �F   ��8�B0���   j j j Q�҃�(��t'_�F    �   ^]� �~ t��P����_^]� _3�^]� ���U���8�H���  ]��������������U���8�H0���   ]��������������U���8�H0�U�E��VWRP���   �U�R�Ћ�8�Q�u���BV�Ћ�8�Q�BVW�Ћ�8�Q�J�E�P�у�_��^��]������������U���8�H0���   ]��������������U���8�H0���   ]��������������U��Ej0P������]��������������U��Ej0P�B�����P������]�����U��E�M��j0PQ�U�R�G�����P�^�����8�H�A�U�R�Ѓ���]�������U��E�M�U��j0PQR�E�P�s�����P������8�Q�J�E�P�у���]��U��Ej$P�����3Ƀ�������]����U��Ej$P������P�����3Ƀ�������]�����������U��E�M��Vj$PQ�U�R�v�����P������83Ƀ��B�P����M�Q�҃���^��]��������U��E�M�U��Vj$PQR�E�P������P�9�����83Ƀ��B�P����M�Q�҃���^��]����U���8�H�U�E���   RPj �у�]���������������U���8�H�U�ER�UP���   Rj �Ѓ�]�����������U���8�P4�E�I�R,P�EP�EPQ�҃�]� ���������U���8�P4�E�I�R0P�EPQ�҃�]� ������������̡�8�P4�A�J4P��Y��������������U��U��V��EP�M�QR���d�����8�H0�E�P� R�U�R�U�R�U�R�U�R�VP�AhR�Ѓ��} ^t(�} t(�E�M�;�~<�U��;�}3�E�M�;�~)�U���} u�E�M�;�~�U��;�}�   ��]� 3���]� �����������U��E��SVW��u�Y��8�P�}���   j hdiuM���Ћ���tK;3u	_^3�[]� ��8�Q���   j hIicM����;�u��8�Q���   j h1icM���Шu��3_^�   []� �����U���8�P�BT��(V�uhfnic���Ѕ�t��8�Q�ȋ��   j
�Ѕ���   ��8�Q�RPhfnic�E�P����P�M������M�藱���u�E�P��虱���M�聱����8�Q�B ���Ѓ��t��8�Q�B ���Ѕ�u��8�Q�B$hfnic���Ћ�8�E�Q�R8Pj
����^��]���������U���8�P0�E�IP�EP�EP�EPQ���   �у�]� ��U���8�P0�E�IV�p� ���   V�uj j j V�uVj Pj=Q�҃�(^]� ����U���8�P0�E�IV�p� ���   V�uV�uj j j�Vj Pj=Q�҃�(^]� ���̡�8�I�P0���   j j j j j j j j j6Q�Ѓ�(�������U��V���4,��8�H0�WVh '�ҋ}�F�E�F    �F   �-�F��8�Q���   ��j hmyal���Ѓ��Ft��t�F    ��8�Q���   j
hhfed���ЉF_��^]� �����������U���8�P�B VW�}�����=ytsdt�MQW������_^]� ��8�B0�N���   Q�ҋ�P������_�   ^]� ��3���������������3�������������������������������3���������������3���������������3���������������3�� �����������U��V���PD�҅�t�E9Ft�F��PH����^]� �����̋A������������̋A��uË ��������������������̸p-�����������U���E�Y(]� ���U���(V���P(�M�Q���ҋN��t&��8�R0j j j j j j P���   j jQ�Ѓ�(��8�Q�J�E�P�ы�8�B�P�M�Q�ҋF����t ��8�Q0�RHj �M�Qj jj?j P�҃���8�H�A�U�WR�Ћ�8�Q�J�E�P�ыF����u3��;��8�E�    �J0�U�Rj j j h  
 j�U�Rh�  jP���   �Ћ}���(��8�Q�J�E�P�у���_u3�^��]Ë�8�B�P�M�Q�ҋF����t ��8�Q0�RHj �M�Qj j j8j P�҃���8�H�A�U�R�ЋF����t��8�Q0jP�BP�Ѓ���8�Q�J�E�P�у��M��I���Ph   h  K j;�U�Rh	��h�  ��跶����8�H�A�U�R�Ѓ��M��k����F��t��8�Q0P�BX�Ѓ��F��t��8�Q0P�BX�Ѓ��F��t'��8�Q0j j j j j jj j jP���   �Ѓ�(j�v$�������   ^��]�����U���SV��W�~j��詃  ��V�^(3ۉ^4�^8�^<��8�H0�Ah�   R�Ћ�8�Q�J�E�P�ы�8�B�PSj��M�h�-Q�҃�SS�E�P�M�Q���E��  �]��i�����8�B�P�M�Q�҃�Sj����  _^[��]���̍A�������������U��VW��~4 tA�I ��8�H��0  h�,hj  ��j
�o�����8�HP�V �AR�Ѓ���uQ9F4u�8�QP�Bh�~0���Ѓ~4 t;��8�Q��0  h�,h�  �Ћ�8�QP�Bl�������m���_3�^]� �M�U�N8�V4��8�PP�Bl�~0���Ѓ~4 t%j
�������8�QP�F �JP�у���u�9F4uۋ�8�BP�PhS���ҋ^<�F<    ��8�PP�Bl���Ћ�[_^]� ��U���8�P�B ��@VW�}�����=MicMtI=fnic��   j�M�蘩���uP���ݩ���M��ũ����8�Q�B4jj����_�   ^��]� ��8�Q���   j hIicM����=�����   htats�M��2�����8�Q�B0j j�M��ЍM�Q�U�R�E�P���E��  �E�    �̴����8���   �
�E�P�у��M������F���F   t��8�J0�QP�҃��EPW���a���_^��]� ���������U��E��V��t3�^]� j�N葀  j�J����F    �v����t��8�H0�QV�҃��   ^]� ��������������j���F�  j�������3�����������U��E3�h�����h  ���P�Ej ��R�Uj PR�s���]� ���������������U��Q�Q��u3���]� �E�H� V�5�8Q�M�Q�E�    �v0PR�V8�ҋ�����t@�E���t9��8�Q�M�RQP�ҋE�����t��8�QW��P�B��W������_��^��]� ������U���8��V��H�A�U�R�ЋU���M�QR���D�������u��8�H�A�U�R�Ѓ�3�^��]� �M�Q�M�L����8�B�P�M�Q�҃���^��]� �������U���8��V��H�A�U�R�ЋU���M�QR��������M���8�P�R8�E�PQ�M�ҡ�8�H�A�U�R�Ѓ���^��]� �������������U���V��M��_I���M�E�PQ���������8���B�U�@<�M�Q�MR�ЍM��J����^��]� ����U���8�P�E���   Vj ��MP��h���h  �j j jj P�EP���S���^]� ��������������U���8V�uW�����   �QV�҃���Vu,��8���   �Q@�ҋ�8�Q4�J P�GP�у�_^]� ��8���   �H�у���u.��8���   �H8V�ы�8�J4�WP�A$R�Ѓ�_^]� ��8�Q��0  h�,h	  �Ѓ�_^]� �����U���4��8�H�QSVW�}W�ҡ�8�P�u���   ��3�SS�Ή]�Ћ�8�QS�E����   j���Ћ�;��M  �d$ �} ~l��8�Q�J�E�P�ы�8�B�Pj j��M�h�-Q�ҡ�8�P�B<�����Ћ�8�Q�RLj�j��M�QP���ҡ�8�H�A�U�R�Ѓ���8�Q0�E����   VP�M�Q�ҋ��8�H�A�U�R�Ћ�8�Q�J�E�PV�ы�8�B�P�M�Q�ҡ�8�P�B<�����Ћ�8�Q�RLj�j��M�QP���ҡ�8�H�A�U�R�Ћ�8�Q�u���   �E��j ��
S���Ћ�8�Q���   �E�j �CP���ҋ����������_^[��]���������������U��E�PV��3Ƀ8������t�   3�h�����h  ���Pj ��Qj R�UR���{���^]� ������U��E3҃8�@V�u ��V�uVR�UR�UR�UR�UPR�?���^]� ����������U��E�E43҃8��R�U<R�U(���\$�E,�$R�E �� �\$�E�\$�E�\$�@�E�$P�2���]�8 ��������������U��E�@3҃8��E��Rj ���T$�$htemf�E �� �\$�E�\$�E�\$�$P�ױ��]�  ���U��E�E 3҃8��R�� �\$�E�\$�E�\$�@�E�$P�Z���]�  ������U��E�@3҃8��E��Rj ���T$�$htcpf�E �� ��'�����\$�E���\$�}�\$�$P�;���]�  �������U��E3҃8��R�UR�UR�UR�UP�EPR����]� U��E3҃8V�u��V��RP�EP�O���^]� ����������U��Q��u3�]� �E�E�H� V�5�8�v0Q�M Q�M���\$���E�$QPR�V(�҃�$^]� ���U���8�P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U���8�P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U���8��P�E���   V���$��MP�ҋ���u�^�    ^]� ��u�^����D{�   ^]� ��^]� ������U���0���8�U�V�U���M�]�P���   �E�PQ�M�E�P�ҋ���̉�P�Q�P�Q�P�Q�P�@�Q�A����  ^��]� ��������U��� ���8�]�V���M�]��P���   �E�PQ�M�E�P�ҋ���̉�P�Q�P�@�Q�A����  ^��]� �����U���VW�};}�M�us��8�P�u���   j htsem���Ѕ�uS��8�QP���   hrdem���Ѕ�u6�MQ�M�U�R�E�}�E�������t�E�M�P�w  _�   ^��]� _3�^��]� U���VW�};}�M�us��8�P�u���   j htsem���Ѕ�uS��8�QP���   hrdem���Ѕ�u6�MQ�M�U�R�E�}�E��ײ����t�E�M�P��  _�   ^��]� _3�^��]� U���SVW�};}��uz��8�P�u���   j htsem���Ѕ�uZ��8�QP���   hrdem���Ѕ�u=��M�Q�]��M�U�R�}��E�腲����t�E������$�  _^�   [��]� _^3�[��]� ��������U���4�ESW�};ǉM�t;Et	;E��   ��8�P�]���   j htsem���Ѕ���   ��8�QP���   hrdem���Ѕ�uj�M��U�U܉E��UԉE��]̉E�M�E�P�M�Q�M�U�U�R�E�P�}�������t+�E̋M�������E��X�E��X��  �   _[��]� _3�[��]� ��������U���SVW�};}����   ��8�P�u���   j htsem���Ѕ�uj��8�QP���   hrdem���Ѕ�uM��U�M��]���Q�M�]��E�R�E�P�}��h�����t%�E��������E��X�  �   _^[��]� _^3�[��]� ���̋A���X(Q�ȋB$��j j h����������������������U���8��0VW���H�A�U�R�Ћ�8�Q�J�E�P�ыE���U�RP�M�Q�M�,�����8�J�U�RP�A�Ћ�8�Q�J�E�P�ы�8�B�P�M�Q�ҡ�8�H�Q��V�ҡ�8�H�A�U�VR�Ѓ�����  ��8�Q�J�E�P�у�_^��]� ������������U���SVW�};}����   ��8�P�u���   j htsem���Ѕ�ue��8�QP���   hrdem���Ѕ�uH��8�Q�J�E�P�ыM���U�R�E�P�}��E�    �-�����u ��8�Q�J�E�P�у�3�_^[��]� ���U��R蛊�����  ��8�H�A�U�R�Ѓ�_^�   [��]� ��U��V�u���  ��^]� �����������U���L��8SV��H�A�U�R�Ћ�8�Q�J3�Sj��E�h�#P���F(��'��S�U�SR�E��  �]�� P�E�P������P�M�Q�1�����P�U�R���R�����8�H�A�U�R�Ћ�8�Q�J�E�P�ы�8�B�P�M�Q�҃�htats�M��͘����8�P�B0jj�M����F(��8�Q�B,���$j�M��ЍM�Q�U�R�E�P���E��  �]��P�����8���   �
�E�P�у�9^4t^��8�BP�PhW�~0���ҋF4;�t�N8Q�Ѓ��F<�^8�^4���8�B��0  h�,h�  �у���8�BP�Pl����_�M��>���^[��]� ������U�����u�E�    �A]� ��u�Q;Ut�   ]� U�����u�E�    �Y]� ��u�E�Y����D{�   ]� �����������U�����u�E�    �Y�E�Y�E�Y]� ��u-�E�Y����Dz�E�Y����Dz�E�Y����D{�   ]� �����U��V�����u#�E�M�U�F�E�N�V�    �F^]� ��u�MQ�VR��������t�   ^]� �������������U��V��F���4,t��8�Q0P�B�Ѓ��E�F    t	V���������^]� ��������������U��V��~ ��,u��8�H4�V�R�Ѓ��E�F    �F    t	V��������^]� �������U���V��3ɍF��H�������8�M��M����   �RQ�M�QP�ҡ�8���   ��U�R�Ѓ���^��]��������������U��V�����u �    ��8�H�A���UVR�Ѓ��#��u��8�Q�Rx�EP�N�҅�t�   ��8�H�A�UR�Ѓ�^]� �������h9Ph�f ��  ���������������U��Vh9h�   h�f ���  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh9h�   h�f ���f  ����t���   ��t�M�UQR����^]� ���^]� ������������U��Vh9h�   h�f ���  ����t���   ��t�MQ����^]� 3�^]� �Vh9h�   h�f ����  ����t���   ��t��^��3�^����������������U��Vh9h�   h�f ���  ����t���   ��t�MQ����^]� 3�^]� �U��Vh9h�   h�f ���V  ����t���   ��t�M�UQR����^]� ����U��Vh9h�   h�f ���  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh9h�   h�f ����  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh9h�   h�f ���v  ����t���   ��t�MQ����^]� 3�^]� �U��Vh9h�   h�f ���6  ����t���   ��t�MQ����^]� 3�^]� �U��Vh9h�   h�f ����  ����t���   ��t�M�UQR����^]� 3�^]� �������������Vh9h�   h�f ���  ����t���   ��t��^��3�^����������������U��Vh9h�   h�f ���f  ����t���   ��t�MQ����^]� 3�^]� �U��V�u�> t3h9h�   h�f �   ����t���   ��t�Q�Ѓ��    ^]���������������U���8�H �Ah]�����������������U���8�H@�AV�u�R�Ѓ��    ^]�������������̡�8�H �������U��V�u���t��8�Q P�B�Ѓ��    ^]���������U���8�P �EPQ�J4�у�]� ����U���8�P �EPQ�J�у�]� ����U���8�P �EPQ�J�у�]� ���̡�8�P �BQ��Y�U��V�uW����������8�H �QVW�҃�_��^]� �����U���8�P �EPQ�J �у�]� ���̡�8�P �B,Q�Ѓ���������������̡�8�P �B0Q�Ѓ����������������h9Ph���P  ���������������U��h9jh���,  ����t
�@��t]��3�]��������U��h9jh����  ����t
�@��t]��3�]��������U��E��u]ËU��� R�UR�UR�UR��]�����������U��E��u��8�H�]Ë��B]��U��E��u]Ë��P]�����������̋�� �-�@�@А�@ ��@ �����������������U��EVh9��jh���F�#  ����t�@��t�M��VQ�Ѓ�^]� 3�^]� �����������̃��� ���������̡�8�H�������3���������������U���8���   �BXQ�Ѓ���u]� ��8�Q|�M�RQ�MQP�҃�]� ���U���8���   �BXQ�Ѓ���u]� ��8�Q|�M�R8Q�MQP�҃�]� ���U��EV��j ���8�Qj j P�B�ЉF����^]� ��̡�8Vj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� ��8�Q�MP�EP�Q�JP�у��F�   ^]� ���̡�8�H���   ��U���8�H���   V�u�R�Ѓ��    ^]����������̡�8�P���   Q�Ѓ�������������U���8�P�EPQ���   �у�]� ̡�8�H�������U���8�H�AV�u�R�Ѓ��    ^]��������������U���8�H�AV�u�R�Ѓ��    ^]��������������U���8�P��Vh�  Q���   �E�P�ы�8���   �Q8P�ҋ��8���   ��U�R�Ѓ���^��]��������������̡�8�P�BQ�Ѓ����������������U���8�P�EPQ�J\�у�]� ����U���8�P�EP�EP�EP�EP�EPQ���   �у�]� �U���8�P�EP�EP�EP�EPQ�JX�у�]� �������̡�8�P�B Q��Y�U���8�P�EP�EP�EP�EPQ���   �у�]� �����U���8�P�EP�EP�EPQ�J�у�]� ������������U���8�H��   ]��������������U���8�P�R$]�����������������U���8�P��x  ]��������������U���8�P�EP�EP�EP�EPQ�J(�у�]� ��������U���8�P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U���8�P�EP�EP�EP�EPQ�J,�у�]� ��������U���8V��H�QWV�ҋ���8�H�QV�ҋ�8�Q�M�R4Q�MQ�MQ���W���Pj j V�҃�(_^]� �����������U���8�P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U���8�P�EP�EPQ�J@�у�]� U���8�P�EPQ�JD�у�]� ���̡�8�P�BLQ�Ѓ���������������̡�8�P�BLQ�Ѓ���������������̡�8�P�BPQ�Ѓ����������������U���8�P�EPQ�JT�у�]� ����U���8�P�EPQ�JT�у�]� ����U���8�P�EP�EPQ���   �у�]� �������������U���8�P�E���   ��VP�EPQ�M�Q�ҋu�    �F    ��8���   j P�BV�Ћ�8���   �
�E�P�у� ��^��]� ������̡�8�P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡�8�H�������U���8�H�AV�u�R�Ѓ��    ^]��������������U���8�P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U���8�P�EPQ�J�у�]� ���̡�8�P�BQ��Y�U���8�P�EP�EPQ�J�у�]� U��VW���t����M�U�x@�EPQR���^����H ���_^]� �U��VW���D����M�U�xD�EPQR���.����H ���_^]� �V�������xH u3�^�W�������΍xH������H �_^�����U��V�������xL u3�^]� W���Я���M�U�xL�EPQR��躯���H ���_^]� �������������U��V��蕯���xP u���^]� W�������M�U�xP�EP�EQRP���e����H ���_^]� ��������U��V���E����xT u���^]� W���/����M�xT�EPQ�������H ���_^]� U���S�]��VW��t.�M�膄���������xL�E�P�������H ��ҍM�������}��tZ��8�H�A�U�R�Ћ�8�Q�J�E�WP�ы�8�B�P�M�Q�҃���艮���@@��t��8�QWP�B�Ѓ�_^[��]� ������U��V���U����x` u
� }  ^]� W���=����x`�EP���/����H ���_^]� ��U��VW�������xH�EP�������H ���_^]� ���������U��SVW�������x` u� }  �#���ϭ���x`�E���P��輭���H ��ҋ���8�H�]�QS�҃�;�A��8�H�QS�҃�;�,�������M�U�xD�EPQSR���h����H ���_^[]� _^�����[]� ��������������U��V���5����xP u
�����^]� W�������M�U�xP�EP�EQ�MR�UPQR��������H ���_^]� ��������������U��V���լ���xT u
�����^]� W��转���M�xT�EPQ��諬���H ���_^]� ��������������U��V��腬���xX tW���w����xX�EP���i����H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u��]  ����t.�E�;�t'��8�J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡�8�H��   ��U���8�H��$  V�u�R�Ѓ��    ^]�����������U���8�UV��H��(  VR�Ѓ���^]� �����������U���8�P�EQ��,  P�у�]� �U���8�P�EQ��,  P�у������]� ���������̡�8�H��0  ���8�H��4  ���8�H��p  ���8�H��t  ��U��E��t�@�3���8�RP��8  Q�Ѓ�]� �����U���8�P�EPQ��<  �у�]� �U���8�P�EP�EP�EPQ��@  �у�]� ���������U���8�P�EP�EPQ��D  �у�]� �������������U���8�P�EPQ��H  �у�]� �U���8�P�E��L  ��VWPQ�M�Q�ҋu����8�H�QV�ҡ�8�H�QVW�ҡ�8�H�A�U�R�Ѓ�_��^��]� ��������������̡�8�P��T  Q�Ѓ�������������U���8�P�EPQ��l  �у�]� ̡�8�P��P  Q�Ѓ�������������U���8�P�EPQ��X  �у�]� ̡�8�H��\  ��U���8�H��`  V�u�R�Ѓ��    ^]�����������U���8�P�EP�EP�EP�EP�EPQ��d  �у�]� �U���8�P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���w���2!����3��F�F �F$�F(�F,�F0�F4�F8�F<�F@�FD�FH�FL�FP�FT�FX�_p��G`�Gd�Gh�Gx�����G|   ��_^��������������V��W�>��t7��������xP t$S������j j �XPj�FP���ݧ���H ���[�    �~` t��8�H�V`�AR�Ѓ��F`    _^������������U��SV��Fx��8�Q��   WV�^dSP�EP�~`W�у����F|��   �> ��   �; ��   �U�~pW�^hSR�Լ������u#���h�-��8�H��0  h�   �҃��E�~P����#���j j jW�^������F|t��������F|_^[]� �F|_�Fx����^[]� �F|�����    ��8�Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��V��~d �F`tLW�};~xtBWPj�NQ��������F|u�E���~xt�    �F`_^]� �M���Fx����t�3�_^]� U��QVW�}�����Y  ��8�H�QhV�҃�����8u"�H��0  h�-h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���t�3�9u�~!�E���<� t��Q����W  �E��;u�|�UR�+�����_�   ^��]� �����������U��QVW�}����>Y  ��8�H�QhV�҃�����8u"�H��0  h�-h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���tЋE��t�3�9u�~:��E�<� t'����8�QP�Bh�Ѓ���t�M��R����V  ��;u�|ȍEP�K�����_�   ^��]� �����������h�-h�   hD�h�   ��������t�������3��������V���(����N^�������������������U��VW�}�7��t��������N���V��������    _^]�U��E�M�UP��P�EjP胹����]��������������̸   �����������U��V�u��t���u8�EjP脹������u3�^]Ë��q�����t���t��U3�;P����#�^]�����h9Ph^� �������������������U��Vh9jh^� ���y�������t�@��t�M�UQRV�Ѓ�^]� 3�^]� �Vh9jh^� ���<�������t�@��tV�Ѓ�^�3�^���U��Vh9jh^� ���	�������t�@��t�M�UQRV�Ѓ�^]� ���^]� U���  Vh9jh^� �����������t/�@��t(�MWQ��x���VR�Ћ��E���b   ���_^��]� �u���x���N`�x�����   � x����   ��w����ݞ�  ��^��]� ����U��Vh9jh^� ���9�������t�@��t�M�UQRV�Ѓ�^]� ��������U��Vh9jh^� �����������t�@��t�M�UQ�MRQV�Ѓ�^]� ����U��Vh9j h^� ����������t�@ ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh9j$h^� ���i�������t�@$��t�MQV�Ѓ�^]� 3�^]� �����U��Vh9j(h^� ���)�������t�@(��t�M�UQ�MR�UQRV�Ѓ�^]� U��QVh9j,h^� �����������t �@,���E�t�E�MPQV�U���^��]� ��^��]� ��������U��Vh9j0h^� ����������t#�@0��t�E�M�U���$QRV�Ѓ�^]� 3�^]� ��������Vh9j4h^� ���L�������t�@4��tV�Ѓ�^�3�^���Vh9j8h^� ����������t�@8��tV�Ѓ�^�������U���`Vh9jDh^� �����������t(�@D��t!W�M�VQ�Ћ��E���   ���_^��]� �u���=u����^��]� ����U��Vh9jHh^� ����������t�@H��t
�MQV�Ѓ�^]� ������������U��Vh9jLh^� ���I�������t�@L��t�MQV�Ѓ�^]� ���^]� ����U��Vh9jPh^� ���	�������t�@P��t
�MQV�Ѓ�^]� ������������U��Vh9jTh^� �����������t�@T��t
�MQV�Ѓ�^]� ������������U��Vh9jXh^� ����������t.�@X��t'�M �UQ�MR�UQ�MR�UQ�MRQV�Ѓ� ^]� 3�^]� �������������Vh9j`h^� ���,�������t�@`��tV�Ѓ�^�3�^���U��Vh9jdh^� �����������t�@d��t�MQV�Ѓ�^]� 3�^]� �����U���Vh9jhh^� ����������t1�@h��t*�MQ�U�VR�Ћu��P�������M��������^��]� �u��������^��]� �����������Vh9jph^� ���L�������t�@p��tV�Ѓ�^Ã��^��Vh9jlh^� ����������t�@l��tV�Ѓ�^Ã��^��Vh9jth^� �����������t�@t��tV�Ѓ�^�3�^���U��Vh9jxh^� ����������t�@x��t
�MQV�Ѓ�^]� ������������Vh9j|h^� ���|�������t�@|��tV�Ѓ�^�������Vh9h�   h^� ���I�������t���   ��tV�Ѓ�^�U��Vh9h�   h^� ����������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������U��Vh9h�   h^� �����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U���Vh9h�   h^� ���s�������tU���   ��tKW�M�VQ�Ћ�8�u���B�HV�ы�8�B�HVW�ы�8�B�P�M�Q�҃�_��^��]� ��8�H�u�QV�҃���^��]� ����������Vh9h�   h^� �����������t���   ��tV�Ѓ�^Ã��^������������U��Vh9h�   h^� ����������t���   ��t
�MQV�Ѓ�^]� ������U��Vh9h�   h^� ���V�������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh9h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������Vh9h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������U��Vh9h�   h^� ���v�������t%���   ��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���U��Vh9h�   h^� ���&�������t���   ��t�M�UQRV�Ѓ�^]� ���^]� ����������U��Vh9h�   h^� �����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh9h�   h^� ����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh9h�   h^� ���6�������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh9h�   h^� �����������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������Vh9h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������Vh9h�   h^� ���Y�������t���   ��tV�Ѓ�^�3�^�������������Vh9h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������Vh9h�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������U��Vh9h�   h^� ����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������Vh9h�   h^� ���I�������t���   ��tV�Ѓ�^�3�^�������������U���Vh9h�   h^� ����������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh9h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ��Vh9h�   h^� ���I�������t���   ��tV�Ѓ�^�3�^�������������U���Vh9h�   h^� ����������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh9h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ��Vh9h�   h^� ���I�������t���   ��tV�Ѓ�^�3�^�������������U��Vh9h�   h^� ����������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��QVh9h�   h^� ����������t#���   ���E�t�E�MPQV�U���^��]� ��^��]� ��U��Vh9h�   h^� ���f�������t!���   ��t�E�M�U���$QRV�Ѓ�^]� ���������U��Vh9h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh9h�   h^� �����������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh9h   h^� ���v�������t��   ��t�MQV�Ѓ�^]� 3�^]� ���������������Vh9h  h^� ���)�������t��  ��tV�Ѓ�^�3�^�������������U���Vh9h  h^� �����������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh9h  h^� ���c�������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh9h  h^� �����������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U��Vh9h  h^� ���f�������t��  ��t
�MQV�Ѓ�^]� ������U��Vh9h  h^� ���&�������t��  ��t
�MQV�Ѓ�^]� ������U��Vh9h  h^� �����������t��  ��t
�MQV�Ѓ�^]� ������Vh9h   h^� ����������t��   ��tV�Ѓ�^�3�^�������������U��Vh9h$  h^� ���f�������t��$  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh9h(  h^� ����������t!��(  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh9h,  h^� �����������t��,  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh9h0  h^� ���y�������t��0  ��tV�Ѓ�^�3�^�������������U��Vh9h4  h^� ���6�������t��4  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh9h8  h^� �����������t��8  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh9h<  h^� ����������t��<  ��t�M�UQ�MRQV�Ѓ�^]� ��������������U��Vh9h@  h^� ���F�������t��@  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh9hD  h^� �����������t��D  ��tV�Ѓ�^�3�^�������������U��Vh9hH  h^� ����������t��H  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh9hL  h^� ���f�������t��L  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh9hP  h^� ����������t!��P  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��QVh9hT  h^� �����������t'��T  ���E�t�E�M�UPQRV�U���^��]� ��^��]� ��������������U��Vh9hX  h^� ���f�������t%��X  ��t�E�M�U���$Q�MRQV�Ѓ�^]� �����U��Vh9j<h^� ����������t�@<��t�M�UQRV�Ѓ�^]� ��������U��Vh9j@h^� �����������t�@@��t�MQV�Ѓ�^]� 3�^]� �����h9Ph�� �������������������h9jh�� ��������uË@����U��V�u�> t/h9jh�� �S�������t��U�M�@R�Ѓ��    ^]���U��Vh9jh�� ����������t �@��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh9jh�� �����������t�@��t�M�UQR����^]� ����������U��Vh9jh�� ����������t�@��t�M�UQR����^]� ����������U��Vh9jh�� ���I�������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh9j h�� �����������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh9j$h�� ����������t �@$��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh9j(h�� ���Y�������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh9j,h�� ���	�������t0�@,��t)�M$�E�UQ�M���\$�E�$R�UQR����^]�  3�^]�  �����������U��Vh9j0h�� ����������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh9j4h�� ���Y�������t5�@4��t.�M(�E �UQ�M���$R�UQ�MR�UQ�MRQ����^]�$ 3�^]�$ ������U��QVh9j8h�� �����������t�@8���E�t�E�MPQ���U�^��]� ��^��]� ����������U��Vh9j<h�� ����������t�@<��t�M�UQR����^]� ����������U��Vh9j@h�� ���i�������t�@@��t�M�UQR����^]� 3�^]� ���U��Vh9jHh�� ���)�������t�@H��t�M�UQR����^]� 3�^]� ���U��Vh9jDh�� �����������t�@D��t�M�UQR����^]� 3�^]� ���U��QVh9jLh�� ����������t#�@L���E�t�E�EP�����$�U�^��]� ��^��]� �����U��Vh9jPh�� ���Y�������t�@P��t�M�UQR����^]� 3�^]� ���U��Vh9jTh�� ����������t �@T��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh9jXh�� �����������t(�@X��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh9j\h�� ���y�������t(�@\��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��V��~ Wu h9jh�� �"�������t�@�ЉF�~��t6h9jh�� ���������t�@��t�M�UVQ�MRQ����_^]� _3�^]� ��������������U��V��W�~��t+h9jh�� ��������t�@��t�M�UQR���Ѓ~ t1h9jh�� �p�������t�N�U�M�@R�Ѓ��F    _^]� ����������U��V��~ u h9jh�� �#�������t�@�ЉF�v��t+h9jh�� ���������t�@��t�M�UQR����^]� �������������U��V�q��t@h9jh�� ��������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ��������������U��V�q��t<h9j h�� �T�������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U��SV��~ Wu h9jh�� ��������t�@�ЉF�}�]�M�UWSQR���<  ��t�N��t�E�UWSPR����_^[]� _^3�[]� �U��V�q��t8h9j(h�� ��������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� ������U��I��t)�E$�E�UP�E���\$�E�$R�UPR����]�  3�]�  �������U��V�q��t<h9j0h�� ��������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U��E��u�E�M�$9� 9�   ]� �����������U��E�����V��   �$���   ^]á(9�����(9uT�EP�3�����=�.  }�����^]Ëu��t�h�-jmhD�j览������t ���������9tV�������   ^]��9    �   ^]ËM�UQR��E������������^]�^]�jE���-(9u.�E���7z���9��t������V�`������9    �   ^]Ã��^]Ð2�����*���������������̡�8�H\�������U���8�H\�AV�u�R�Ѓ��    ^]�������������̡�8�P\�BQ�Ѓ���������������̡�8�P\�BQ�Ѓ����������������U���8�P\�EPQ�J�у�]� ����U���8�P\�EP�EPQ�J�у�]� U���8�P\�EPQ�J�у�]� ���̡�8�P\�BQ�Ѓ����������������U���8�P\�EPQ�J �у�]� ����U���8�P\�EP�EPQ�J$�у�]� U���8�P\�EP�EP�EPQ�J(�у�]� ������������U���8�P\�EPQ�J0�у�]� ����U���8�P\�EPQ�J@�у�]� ����U���8�P\�EPQ�JD�у�]� ����U���8�P\�EPQ�JH�у�]� ���̡�8�P\�B4Q�Ѓ����������������U���8�P\�EP�EPQ�J8�у�]� U���8�P\�EPQ�J<�у�]� ����U���SVW�}��j �ωu������8�H\�QV�҃���S�����3���~?��I ��8�H\�U�R�U��EP�A(VR�ЋM��Q���h���U�R���]����;�|�_^[��]� �������������U���VW�}�E��P������}� ��   ��8�Q\�BV�Ѓ��M�Q������E���taS3ۅ�~L�I �UR���e���E�P���Z���E;E�#����8�Q\P�BV�ЋE����;E��E~߃�;]�|�[_�   ^��]� _�   ^��]� ������������U��M�EV�u������t#W���    �Pf�y������f�8f�u�_^]� �U��� �E���M��"  �ȉES���V�u��W�}�ǃ��Q���ƃ��։E��B��E���؉M�E��U���M��~�U�U���)}�M��>���E��}�t�u+���I �\�P���m���u�E�����E��   )}��u��	;]��u��s���u;]�]�}�M��>P�E�V�Ѕ�}	�u���]�M��E��VP�҅��V������F��}�t!�M�+ȃ����\�P���m���u�]��;]~�����_^[��]� ���U���(W�}�����E�E���M��  �MS�؉E������ǃ��S�����E�ы���V�]�U��E܉U���]��~�E�E��)}��]��)�M�U��E�Q�M�RP������E�����E��   )}��u�;E��؉u�s���u;]�]�}�M���>P�E؋V�Ѕ�}	�u؃��]��M���E�VP�҅��i����}���F�t&�M�+ȃ���I �Pf�\����f�f�u�]��}�;E�w����%���^[_��]� ��������U���(W�}�����E�E���M��)  �ЉE������ǃ��J���SV�uƃ��ΉE��A��E����؉U��E܉M����I �U���~�M�M��)}��U��A�M�ɋE��M�t�M�+���I �\�p���m���4u�E�����E��   )}��u�;E��؉u�s���u;]�]�}�M��>P�E؋V�Ѕ�}	�u؃��]��M��E�VP�҅��Q����}���F�t�M�+ȃ���\�P������u�]��}�;E~�����^[_��]� ���������������U��E�Pu�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����E��SV��W�]�t8�u��t1�}��t*�} t$�VP��Ѕ���   |������E�   �}}_^3�[��]� �}�M���E�������uu��VP�҅�t#}����}����}��E9E�~�_^3�[��]� ��~3�E���]��]�E��E�M���؋ESP���҅�u�����_��^[��]� ���������������U����E��SV��W�]��  �u����   �}����   �} ��   �VP��Ѕ���   }�M_^�    3�[��]� �O�3����E�   �M} ����   �E���8_^3�[��]� ���M�U���<�M������uuVQ���҅�t}�O��M��W�U��M9M�~�뤅�~3�E���]��]�E��E�M���؋ESP���҅�u�����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� �����������U��M�A8��   �IXV�AP�I@���I�AP�I(�AX�I ���I0���A@�I �A8�I(���IH����������Dz�u�؋��eJ����^��]���W���A�IX�AP�I�A8�I�A�I@�AP�I@�U��A8�IX�]������IH�����I0�����e��	����ݝx����A�I(�U��A�I �U��AX�I �]��AP�I(�����IH�E����	���������I�������]��A8�I(�A@�I �����	�������I���E��e��I0�������]��E��e����]����e��ˋE��x������]������]��AH�I@�A0�IX�����]��AX�I�AH�I(�����]��A0�I(�A@�I�����]��AP�I0�AH�I8�����]��AH�I �AP�I�����]��A8�I�A0�I �   �����]��_^��]�������U��y0 tL��E�A�A �A�A(�A��$����������X�X�A� �A �`�A(�`�E����X�X]� ��E����������P���P�E����X�X]� ��̋�3ɉ�H�H�H�V��V�7w���FP�.w��3����F�F^��3���A�A�A����A�`�
�@�b�	���B�a�������U����   ��UV���q�U�W3��<��M��}���  ��S�]�k  ��؋�U��M�U��U�@�����@�U��@�B�@�������@���@�G�>��w����U���  �w������݃��B��   �U������ɋP��R�э����]��B���B�P���R���U����E������]��E��M��E������������]��E����E����E��E��]����E��]����E��]��]����U��E��U�����B���B���U������������]��E����E����������E������E��E��]����E��]����E��]����U��E��]���R�э�������B���B�P���R���U����E��������]��E����E����������E������E��E��]��E��]����E��]��U��E��]�����B���B���U����E��������]��E����E����������E������E��E��]��E��]����E��]��E��U��`�����E�U���������;���   �ލ�+���͋�@����������]��@���]��@���U������M������]��E��E����E��������]��E������������E��E��]��E��E��]����E��]��E��U�u�������������������������������M���Q�ʍU��R���[�[�+�����E�KH��P�E��SL��H�щKP�P�ST�H�KX�P�������S\z^�E�����������zP���CP�����CX���CH���CX�������cH���[�[ �[(�C(�KP�C �KX���C�KX�C(�KH���CH�K �\���E���������za�CX�����CP�����cH�CH���CP�������[���[ �[(�CP�K(�C �KX���C�KX�CH�K(���C �KH�C�KP�����[0�[8�[@�[�CP�����CX�����KH�CX�����cP���[0�[8�[@�C8�KX�C@�KP���C@�KH�CX�K0���CP�K0�C8�KH�����[�[ �[(��$���SP������E��U�   �����}��M�����م�~�A8����u��1���U�@���K�I��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�@�K@���CX�H�D��@�����U���]��C���@�K0���CH�H���C ��C�@�K8���@�KP���C(��C�C@�H���CX�H3������U��x  �A������܃��E����E   �E�
���������ɋE������׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H�E������������������������������E����]��E��]����]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H�E��������]������M������������������������]��E��]��E��]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H���]������M������������������������]��E�Eȃ��]���E����]ȃE׃m����@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H���]������M������������������������U��E��]��E��U�������E������������;���   �P�U��+ЉU�
���������ʋE���׋��U�@���K��@�K0���CH�H���]�� �K �C�@�K8���@�KP���]�� �K(�C�C@�H���CX�H�   E)E���]����E��������������������M����������]��E��E��U�����[������_��^��]� ��[��_��^���؋�]� �����������h,9Ph_� �������������������h,9jh_� �o�������uË@����U��V�u�> t/h,9jh_� �C�������t��U�M�@R�Ѓ��    ^]���U��Vh,9jh_� ���	�������t�@��t�MQ����^]� 3�^]� �������U��Vh,9jh_� �����������t�@��t�MQ����^]� 3�^]� �������U��Vh,9jh_� ����������t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh,9jh_� ���9�������t�@��t�MQ����^]� 3�^]� �������U��Vh,9j h_� �����������t�@ ��t�MQ����^]� 3�^]� �������U��Vh,9j$h_� ����������t�@$��t�MQ����^]� 2�^]� �������Vh,9j(h_� ���|�������t�@(��t��^��3�^������Vh,9j,h_� ���L�������t�@,��t��^��3�^������U��Vh,9j0h_� ����������t�@0��t�MQ����^]� 3�^]� �������U��Vh,9j4h_� �����������t�@4��t�M�UQR����^]� ���^]� ��Vh,9j8h_� ����������t�@8��t��^��3�^������U��Vh,9j<h_� ���i�������t�@<��t�MQ����^]� ��������������U��Vh,9j@h_� ���)�������t�@@��t�MQ����^]� ��������������U��Vh,9jDh_� �����������t�@D��t�MQ����^]� 3�^]� �������U��Vh,9jHh_� ����������t�@H��t�MQ����^]� ��������������Vh,9jLh_� ���l�������t�@L��t��^��3�^������Vh,9jPh_� ���<�������t�@P��t��^��3�^������Vh,9jTh_� ����������t�@T��t��^��^��������Vh,9jXh_� �����������t�@X��t��^��^��������Vh,9j\h_� ����������t�@\��t��^��^��������U��Vh,9j`h_� ���y�������t�@`��t�M�UQR����^]� 3�^]� ���U��Vh,9jdh_� ���9�������t�@d��t�M�UQR����^]� 3�^]� ���U��Vh,9jhh_� �����������t�@h��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh,9jlh_� ��詿������t�@l��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh,9jph_� ���Y�������t�@p��t�M�UQR����^]� 3�^]� ���U��Vh,9jth_� ����������t�@t��t�M�UQR����^]� 3�^]� ���U��Vh,9jxh_� ���پ������t�@x��t�M�UQR����^]� 3�^]� ���U��Vh,9j|h_� ��虾������t�@|��t�MQ����^]� 3�^]� �������U��Vh,9h�   h_� ���V�������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh,9h�   h_� ����������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh,9h�   h_� ��覽������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh,9h�   h_� ���F�������t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U���|��A�����U����U����U��  S�V�E��EW�����������   ���������U�r�z�
�R;��4v���4��I�$ȍ��F�R�a���F�a�uB�!�]��B�a�U��B�a�U������������]��E����E����������E��������E��G��$ȍ��]��B�a�U��B�a�U������������]��E����E����������E��������E��������m�������_�U�^��[�U����U�������������������蘢 ����������D�Ez���P�P���]� �������E�����E����X�M��X��]� �������U���@��$�A�������E�    ���]����]��]���$�������]����]��]���   �	S�]VW�M��E����������t[��%�����E�M�����@��P�9���F�@��R�M��9���~���Q�M��y9���v;�t�v��P�M��c9���M����m��M�u�_^[�M�UQR�M��A�����]� ����������̋Q3���|�	��t��~�    t������u��3�������U��QV�u;��}�	���    u����;�|���^]� +ƃ�^]� �������U��VW�}��|-�1��t'�Q3���~�΍I �1�������;�t����;�|���_^]� �������������̋Q3���~%V�1�d$ ���   @u�����t������u�^�̋QV3���~�	�d$ ����Шt������u��^�������U��Q3�9A~��I ��$��������;A|�Q��~[SVW�   3ۋ���x5��%���;��E���}$��������%���;E�u�
   ���;q|݋Q���G���;�|�_^[��]�������U��	����%�����E��   @t����������wg�$�h��E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� ��-�A�U�����U����S��V������   @Wt���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V��V�`���FP��_��3����F�F^��U��SV��WV��_���^S��_���E3���;ǉ~�~t_��8�Q���   h(.��jIP�у�;ǉt9�}��t;��8�B���   h(.��    jNQ�҃����uV�k_����_^3�[]� �E�~_�F^�   []� ����������U��SV��WV�2_���^S�)_���}3Ƀ�;��N�N��   9��   �G;���   ��8�Q���  h(.��jlP�у����t=� t@�G��t9��8�Jh(.��    ���  jqR�Ѓ����u���]���_^3�[]� �O�N�G�Q��    R�F�QP�.�������t�N�WP��QPR�.����_^�   []� ���������U��SV��WV�2^���~W�)^��3Ƀ�9M�N�N��   �E;���   ��    ��8�H���  h(.h�   S�҃����t=�} tH�E��tA��8�Q���  h(.��h�   P�у����u���b���_^3�[]� �U�V�,�F   ��8�H���  h(.h�   j�҃����t��E�M�F�PSPQ�-���E����t!�V�?�W�RWP�u-����_^�   []� ��M�_^�   []� ���U��Q2���~CS�]V�1W������������;�u��   @u�����u3���   ��
���u�_^[��]� �����������U��S�]V��3�W�~���F�F�C;CV��   �\��W�~\��3��F�F��8�Q���   h(.jIj�Ѓ������   ��8�Q���   h(.jNj�Ѓ����uV�&\����_��^[]� ��F   �F   ����K�H�C��B�_��^�   []� ��[��W��[��3��F�F��8�B���   h(.jIj�у����t[��8�B���   h(.jNj�у�����\�����F   �F   ����S�Q��K�H��C�B��   _��^[]� �����������U��3�V���F�F�F�EP�������^]� �������������U��EVP���������^]� ����������U���EV���V��������Au��8�H��0  hx.j,�����^��^]� �����U���W������G���U���'������A�  ������A��   ��.������AuR������AuKV��蛣 ��蔣 �ȅ�u��^����__��]Ëƙ����ҋ�u�u��E�^������__��]���������Au������=�.��������Au6�����������U������G�����_��������Au�����U����_�
����������m� �E����U���$��������A{���������__��]�������������__��]����U����.V�E��������At����.������Au�������'����$�$�:� �����'���^�e�����^]� ��������������U����V�E��������u�   �3����]����Az�   �3�3�����$;���W���$����� ��E����$�$謰 �V����������Au��8�H��0  hx.j�����^����_u������������^]� ���U������EV�ы�������z!��8�؋H��0  hx.j5�����U������$�� �]��F�$�� �}��$� � ��E�$�� �^�����&���^��]� ���������������U��M��P]����U��M��P]����U��M��P]����V����.�F    ��8�HP�h��Vhp�h`��҉F����^����������̃y ��.u��8�PP�A�JP��Y��U��A��u]� ��8�QP�M�Rj Q�MQP�҃�]� ��U��A��t��8�QP�M�RQP�҃�]� ������������U��A��t��8�QP�M�RQP�҃�]� �����������̡�8�HP���   ��U���8�HP���   ]�������������̡�8�HP�QP�����U���8�HP�AT]����������������̋��     �@    �V����t)��8�QPP�BL�Ћ�8�QP��J<P�у��    ^�������������U��SV�ً3�;�Wt��8�QPP�B<�Ѓ��3�s�}�Eh��W�C��8�QP�J8hp�h`�P�EP�у�9u�~O�I ���z u!���@   ��8�QP���H�RQ�҃���8�HP��A@VR�Ћ�����;u�A|�3�9_^��[]� ������U��SVW��3�9w~>�]��8�HP��A@VR�Ѓ���t/��8�QPj SjP�B�Ѓ���t��;w|�_^�   []� ��8�QP��JLP�у�_^3�[]� ���������̡�8�PP��JDP�у�������������̡�8�PP��JHP��Y��������������̡�8�PP��JLP��Y���������������U��U�E�@R�URP�I���]� �����U��V��~ ��.u��8�HP�V�AR�Ѓ��Et	V�>W������^]� ����h09Ph�f �p������������������U��h09jh�f �L�������t
�@��t]�����]�������U��Vh09jh�f ����������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R�
����E�NP�у�4�M���4�����^]ÍM�'������^]��U��h09jh�f 謪������t
�@��t]��3�]��������U��h09jh�f �|�������t�x t�P]��3�]������V��F��Wu�~��N�ɍ<u�< ��u_3�^á�8�H�F��  h /j8��    RP�у���tщ~�F_�   ^���U��V��F;Fu������u^]� �N�V�E���   F^]� �����������U��V��FW�};�~ ��|�F�M��_�   ^]� _3�^]� })�V;Vu��������t�F�N��    �F9~|׋V;Vu���������t��F�N�U���F_�   ^]� ������U��V��FW�};�~����}3�;Fu������u_^]� �F;�~�N�T������;ǉ�F�M���F_�   ^]� �U��E��|4�Q;�}-���;Q}V�d$ �Q�t������2;A|�^�   ]� 3�]� ������������U��Q3���V~�I�u91t����;�|���^]� �������V��W�~W�P��3����_�F�F^�����A    ��������̋Q�B���|;�}�QV�4���tP�1�����^�3�����������̍Q3��Q�Q�A�Q�A������������W���O�G;�t#��tV�q��t�~ u3���j�҅���u�^�G�G�G�G    �G�G    _�����U��A��3�;�Vt!��t�M���;�t�@��t
�x t��u�3�^]� ��������U��Q�E�P�Q�P�Q�B�A]� �U��E�Q�P�Q�P�Q�B�A]� ̋Q��3�;�t�ʅ�t�I����t
�y t��u�����������U��E�P�Q�H�A�@�H]� ����U��E�P�Q�H�A�A�H]� ���̋Q��t!�A��t�B�A�Q�P�A    �A    ��������V��W�~W�L/�N��3����_�F�F^��������������U���SV�uW���^S�}��N��3���F�F�O�N�W���V9G�E~��I �O���F9F�U�uL��u�~��~��t���< ��t\��8�H���  h /j8��    RP�у���t3�~�}���V��M����E�F��;G�E|�_^�   [��]� _^3�[��]� �������������U��V�u��|'�A;�} �U��|;�};�t�A��W�<��<���_^]� ���������U��EV�u;�}����|,�Q;�}%��|!;�};�t�QW�<�P������tVW����_^]� ����������U��V�q3���W~�Q�}9:t����;�|���P�����_^]� ���������������U����E�Qj�E��ARP�M��E�T/������]� �����U����Q�Ej�E��A�MRPQ�M��E�T/�������]� ̋A��;�t?W3�;�t7V�H;�t	9yt���3��P;�t;�t�J�H�P�Q�x�x;���u�^_������̋Q����.t!�A��t�B�A�Q�P�A    �A    �̋�� \/�@�.�HV3��q�q�P�r�r��.�p�p�p�P�H^������V���\/�����F3�;��F�.t�N;�t�H�F�N�H�V�V�F;��F�.t�N;�t�H�F�N�H�V�V^�U��E�UP�AR�Ѓ�]� ���������U��V��N3�;���.t�F;�t�A�F�N�H�V�V�Et	V�VN������^]� ������������U��V��W�~W�L/��J��3����E��F�Ft	V�N����_��^]� ������U��V��������Et	V��M������^]� ���������������U���8�PH�EPQ���  �у�]� �U���8�P�B4VW�}j��h�  ���ЋMWQ���D  _^]� ��������������U��V���PXW�ҋ}P���gu�����Et�_�   ^]� �M�UPWQR���1  _^]� �����������U��S�]VW��j ���<s���8�  �}uI�~ uC��8�P���   j h�  ���Ѕ�u��8�QP���   h�  ���Ѕ�t	_^3�[]� �M�U�EQ�MRPSWQ����  _^[]� ��������U��EP�A    ������]� �����̸   �A� ������A   � ������U���@S�]��`��VW��u�G   �}  ����   �M3�V�Jr���8�  u4����P�w蔻����8�P�M�B4��jh�  ��_^�C�[��]� �MV�r���8�  u�E�M��RPQ����_^�   [��]� �MV��q���8�  t�MV��q���8��  ��8�P�M�B4jh�  �Љw�  ����  �E�H��BXj	��P�C��3��؃�;މu�t��8�QH���  VS�Ѓ��E��M�;O�f  9w�]  ��8�B�M���   Vh�  �҅�u!��8�P�M���   Vh�  �Ѕ��  ��8�Q�M�B4Vh�  ��;�t
V���������E��G��8���   ���   �Ћ];މE���   ;���   S�7����M���jQ�ˉu��uĉuȉủuЉu؉u������U�E��ˉu��u�u�U�E��]��E�   ������t!��t��t�u���E�   ��E�   ��E�   ��S���M�;�t�N�����BX�M�Q����P�T���M܃�;�t�L����M���h���M���h���M������]�M�U�EQSRP����  _^[��]� �M�����_^�   [��]� �������������̸   � ��������� ������������̃��� ����������� �������������U���8�H�QV�uV�҃���^]� ̸   � ��������3�� ����������̸   @� ��������3��  ����������̸   � ��������U��W�}��u3�_]� ��U�@@VR�Ћ���u^_]� ��8�Q0�F�M���   PQW�ҋF��^_]� U���8�H0�U�AR�Ѓ���t
��ȋj��]� �������3�� ��������������������������̸   � ��������3�� �����������3�� �����������U��E� ����]� �������������̸   � ��������U��E� ����]� ��������������3�� �����������U���8�H���  ]��������������U���8�H���  ]��������������U���8�P�EP�EP�EP�EPQ���   �у�]� �����U���8�E�P�EP�E���\$�E�$PQ���   �у�]� �������������U���8�P�EP�EP�EPQ���   �у�]� ��������̡�8�P���   Q�Ѓ�������������U���8�P�EP�EP�EPQ���   �у�]� ���������U���8�P�EP�EPQ���   �у�]� �������������U���8�H�U�ApR�Ѓ�]� �����U���8�P�EP�EPQ���  �у�]� �������������U���8�P�EP�EPQ���  �у�]� �������������U���8�P�EP�EPQ���  �у�]� �������������U���8�P�EP�EPQ���  �у�]� �������������U����   V�u��u3�^��]�Wh�   ��0���j P�d� ��R���E�P���ҡ�8�P�B<�M��Ѕ��}t0j �M�QW�!,������u��8�B�P�M�Q�҃�_3�^��]ËE�M�Uh�   ��p�����0���P��t����MQWj	��P�����0���ǅ4���PJ�E��u�E���E� �E��u�E���E��N�E�`%ǅx��� ǅ|����u�E���E��u�E���E���E��E���E���E���E��u�E� O�E�O��L����8���B�P�M�Q�҃�_��^��]����������U���   SV�u(3ۅ��]�u��8�H�A�UR�Ѓ�^3�[��]Ë�8�Q�B<W�M3��Ѕ��'  謄�����E�tq�MQ�M�虴��Wh�*�M�����P�M�肴���u�Wj��U�R�E�P��\���Q�_?�%�����P��x���R�5�����P�E�P�(�����P���������E�t�E� �� t�M����蠴����t��x������荴����t��\�������z�����t�M̃���j�����t��8�Q�J�E�P����у���t�M��@����}� t"�U(�E$�M�R�UP�EQ�MRPQ���������U�R蟃������E$�M�UVP�Ej QRP�����������8�Q�J�EP�у���_^[��]����������������U��E�M�UP�EQ�Mj RPQ������]�������������̋�`<����������̋�`L����������̋�`0����������̋�`P����������̋�`$����������̋�`4����������̋�`D����������̋�`T����������̋�`(����������̋�`H����������̋�`����������̃��  3ĉD$�X+S�\$�T$��@�D$�L$W��   ����   �ً���������   �ً�������uq�ً�������ub��u^8D$uX8D$uR�   �H�3ۃ���   �D�D��T$+ш\$�\$�\$�\$
�L$�+Ȉ�D$_[�L$3��z ��À|$@uK3�:�uE�ы�������u6�ы�������u'������u8\$u8\$u8\$u
3��K�f���h<0h(0h�   h0蛙 ����_�D$�D$�D$�D$�D$�D$	�D$
�D$�D$[�L$3��_y ��Ã�u��D�D��T$+ш\$�\$�\$�\$
�L$+Ȉ��D$�L$_[3��y ����������������Q��0S�\$�L$�T$����<@uF��uB������u9������u0�   �H���ux�D�D��T$+эL$� +�� �D$[YÀ�@u��u������u����u3��H�h�0hl0h�   h0�t� �����D$�D$�D$�D$�D$[YÃ�u��D�D��������̃��  3ĉD$�gfff����������+ʃ�	S�D$0�D$1�D$2�D$3�D$4�D$	5�D$
6�D$7�D$8�D$9�-w	�L�O��_�ȸgfff����������+ʃ�	w	�L�O��_�ȸgfff����������+ʃ�	w	�L�O��_V��gfff��������ʍ��+��	w	�D4�G��_�gfff����������+ʃ�	^w	�D�G��_�L$�[3��G �w ����̋��   ���   �89���   �<9���   ���   �ɣ@9�D9t��3�����SW�|$��tM���tG��0tB�H9��t;V��p����t*����I :u�J������u���: u�> t� ��u�^_[�3�_[����́�   �  3ĉ�$�   ��$�   ��$�   ��$�   SV�5H9�D$��$�   3�;�L$�T$�D$t*���L$Q���   R�/Q  ����t�6;�u��;��x  9T9�l  ��  ��"��Ǆ$�   �^fǄ$�   Qf��$�   Ƅ$�   �Ƅ$�   ���$�   Ƅ$�   Ƅ$�   ���$�   ��$�   ��$�   �D$8�	�vf�D$<Pf�t$>�D$@��\$A�\$B�D$C�D$D��T$E�L$F�D$G�D$x�`Gf�D$|�f�t$~Ƅ$�   �Ƅ$�   ���$�   Ƅ$�   Ƅ$�   ���$�   ��$�   ��$�   �D$X��O�f�D$\f�t$^�D$`��\$a�\$b�D$c�D$d��T$e�L$f�D$g�D$�c�f�D$Kf�t$�D$ ��\$!�\$"�D$#�D$$��T$%�L$&�D$'�D$(��f�D$,*>f�t$.�D$0��D$1�\$2�D$3�D$4��T$5�L$6�D$7�D$H��L-f�D$L*>f�t$N�D$P��D$Q�\$R�D$S�D$T��T$U�L$V�D$W�ĈD$t��$�   ��$�   P�L$Q�D$pC�o�f�D$t*�f�D$vF�D$x��D$y��D$z��D${��D$}��D$~*�D$6Ǆ$�   ��
fǄ$�   4MfǄ$�   �KƄ$�   �Ƅ$�   Ƅ$�   Ƅ$�   NƄ$�   rƄ$�   =Ƅ$�   �Ǆ$�   1c_ffǄ$�   f*fǄ$�   �LƄ$�   �Ƅ$�   �Ƅ$�   �Ƅ$�   �Ƅ$�   �Ƅ$�   �Ƅ$�   TƄ$�   �5N  �����n  �T$8R�D$P�N  �����T  �L$xQ�T$R�N  �����  �D$XP�L$Q��M  �����  �T$R�D$P��M  ����u^�Pf[��$�   3��r �Ĵ   ÍL$(Q�T$R�M  ������   �D$HP�L$Q�M  ������   �T$hR�D$P�gM  ����tl��$�   Q�T$R�NM  ����u^�`e[��$�   3��r �Ĵ   Í�$�   P�L$Q�M  �������^%pd[��$�   3���q �Ĵ   �^��P[��$�   3��q �Ĵ   �^��c[��$�   3��q �Ĵ   �^�H>[��$�   3��q �Ĵ   Ë�$�   ��^[3��hq �Ĵ   �������̍A������������̋D$���   ����   �P���   ���   �P�H� �����̸������������̋�� �0�@    �SW���O3�;�t0V��8\9���   ���   ���   u	��Pj��;��u׉_^_[�SU��V�u3ۅ���   W�|$�FWP�K  ����t�ދ��   ��u�_��^][� ���� ��t�V�� ����tߋ��d� ��3�;�t�;�t���   �;uu	�}���   ���   ���   ���   ���   ��Bj���Ћ�_^][� ��^][� ��������������V�q��t/S�\$W����P<���   S���҅�u��Pj���҅���u�_[^� �����W��� u;�L$�A����   �G�A    �G����   �I ���   ���   ��u�_� U�l$V�u��t(S���   �FP��������t��Bj���Ѕۋ�u�[�M��^�E    ��]t��I ���   ���   ��u��G��u�O_� ���    t���$    ���   ���    u񉈴   _� ������̋A��t���$    ���   ���   ��u����������������̋�V3��ҋȅ�t)�T$3���t!��$    ;�t�I��u�^� �   ^� ��^� �̋D$�`/�d/��h/�P�l/�H�P� �����̋D$�Q��Q�P�Q�I�P�H� �̋D$�Q$��Q(�P�Q,�I0�P�H� �̋D$�Q��Q�P�Q�I�P�H� �̋D$�Q��Q�P�Q�I�P�H� �̋D$�Q��Q�P�Q �I$�P�H� ��V�q��W�   t����P���ҋ��   ���u��_^������̋D$� ��������̋���V�ҋ���tu�F��u�,1W�|$Ph1W�C0 h1W�80 ���   ���   ���   �L$ ���L$�D$���   Q�ωT$�D$�a6 h�&W��/ ��_^��� �T$h�0R��/ ��^��� �̋A��t;�t	��R0����� ��������̃�8�  3ĉD$4�D$@SU�l$DV�t$PW��jP�_j S�|$�l$$�D$ �q jP�GXj P��p �L$DVQ�F  �p�P��@�t$D���   ��V�T$D�� ��V�FtjOUS�+� ���D$��tjOP�GXP�� ���GXP�(������; �Gu1h�2hh2h  h0�ԋ ��_^][�L$43��k ��8� S����������D$��   �=P9~lh2hh2h  h0�U� ���   �|$ ty�|$<���+����D$jOPS�D$N �i� jO��QS�� S�x����|$,������'  �D$|���t1h�1hh2h"  h0�� ��_^][�L$43���j ��8� �;Ou6�	Nu0�
_u*�Ou$�bu�ju�eu�cu�tu� t7�X u1h�1hh2h2  h0裊 ��_^][�L$43��j ��8� ��N���ĉ�V�H�N�P�T9   �H����������T9    t1hd1hh2h;  h0�7� ��_^][�L$43��j ��8� V�)F  ����t1h41hh2hA  h0��� ��_^][�L$43���i ��8� �; tZ�5H9��tP���~ uB�NX��t;�Ð�:u��t�P:Qu������u�3��������u�T$�V����|$�6��u��=H9 t�L9��t�8��=H9�L$D�=L9�    _^][3��Ei ��8� �������0�5��������SV�t$W3�������   9��   ��   U�nUh`/�"D  ����tpU���3�����ud���� ��tBV�n� ����t��ȋBW�Ћ���u*h�2h�2h]  h0讈 ��]��_^[� �   ���   �K���   �s]��_^[� �̋D$SW�x����t?V�( t-����  ����t V�w� ��P��������u��Bj���Ћ��   ��u�^_[� �������������S�\$UV��nW3���~�F�<� ��t� ��ȋB0S�Ѓ�;�|�n(3���~$��I �N$�<� ��t� ��ȋB0S�Ѓ�;�|�n83���~'���    �N4�<� ��t� ��ȋB0S�Ѓ�;�|�nh��~#3����    �Nd�9�B0�S�Ё��   ��u�nX��~3��NT�9�B0�S�Ѓ�h��uꋮ�   ��~3����   �9�B0�S�ЁǨ   ��u䍎�   �e� _^][� �������������̀=�9 �u��9�=�9 �!  j ��9��m  j ��k j �Yl j �l j ��l j �[ j ��� j �N j ��F j �xp
 j �1q
 j �q
 j �p
 j ��p
 j �Uq
 j �>	 ��@j �$	 j �	 j �	 j �o	 j ��	 j �A	 j �w
 j �� j �� j � j �% j � j ��
 j �9� j �� j ��
 ��@j �Q�  j �> j �39 j �ܺ
 j 西	 j ��� j � j �`� j �X j �2k j �kk j ��j j ��
 j �֍
 j ��� j �t
 ��@j �� j �gf
 j �@`
 j �0
 j �� j �k� j ��&
 j �]
 j �F� j �� j ���	 j �q� j �z�	 j �	 j �4 j ���	 ��@j 苼	 j �T�	 j �D  j �q	 j �� j �(� j �� j ��� j �#� j �\� j �� ��,��3�V��L$���   �L$��F�P9���   �T$���   ���   ���   ���   ���   ���   ���   �D$R���   �L$PQ��ǆ�      �������      ���^� ������������V����0�"����D$t	V�u*������^� �����������̋D$V��P��0�F    �f�����^� VW�|$��;�t�����W���G���_��^� �����������̋��t���@á���@����������̋��t���x ��á���x �����V��L$�$ 3Ʌ�tf9t���$    ��f�<H u�PQ���=" ��^� ������̋	����t��3�9P��#ы�á��3�9P��#ы�Ë	��+�����#�����������������3���A�A�A�A�A�A�A �A$�A(�A,�������������̃9 u?�y u9�y u3�y u-�y u'�y u!�y u�y  u�y$ u�y( u	�y, u3�ø   ������̃�4�  3ĉD$0V�t$<W������� ��}2j0�D$j P��f ���L$Qj0���	 _^�L$03��b ��4� �R���" ��t �G�OPQ����" ��t��Wj���# �L$8_^3���a ��4� �����������QS3�UV��L$��^�^W�~�nV�] �^�^�^�^ �^$�^(�^,�7" :ÈD$t"�L$W�" :ÈD$t�L$Uj� �D$�L$�d	 =���|�L$��� ��}���_�] �^�^�^�^ �^$�^(�^,�D$_^][Y� ����VW�|$h�3W���$ ���> uO�~ uI�~ uC�~ u=�~ u7�~ u1�~ u+�~  u%�~$ u�~( u�~, uh�3W�# ��_^� ���/# h�&W�# �j Ph�3W�# �N�VQRh�3W�# �F,�N(�V$P�F Q�NR�VP�FQ�NRPQh\3W�V# ��P���# _^� �������V����t4��;��t���~����uP��>  ������^Ë���^Ë���^����������V����t[��;��tP���~��������^�u��t	�x ~� �@    ^�h44h 4jJh4� ������^Ë���^�VW�����t!��;��t���~����u	P�>  ���t$������~-�NQ�=  �p���    �@    V��j P��c ��_^� ����S��V�3��t��;5��u�D$P�q���^[� �>W�|$~>W�\������t�������F;�|����~KW���KVQ�Pg ���{_^[� ;~~,�WRV�e=  ���F��N��+у�R�j Q�	c ���~_^[� �������������SVW�|$����~]�\$��tU�; tPW�0����WSP��f ��������t������x�6�ƅ�t�H���_� ^[� ���H_� ^[� ��������t����8~������_^[� ����t���@    �_^� [� ���@    �_^� [� VW�|$������   S�\$��ty�; tt���t�������@U�P�V�����-������t����ŋPW�SR��e �����t�����x�6�ƅ�t]���@[_� ^� �ŋ@� ][_^� �������̋T$�ҡ��V��t#�: t��W�x�I �����u�+�RP���l���_��^� ����̡��V��L$�ɉt!f�9 t3���    ��f�<A u�QP���} ��^� ������̡��V��L$��� 3Ʌ�tf9t����f�<H u�PQ���= ��^� �������U�l$V��M 9�
  �������t����x �������������^]� ����t����8 ~C�h'
 ��u4�������E ��t��� �M ���^]� ���� �M ���^]� ����E ��t����PSR�������M �������t����Ëх�W�xt�����3�9BW����#�Q�Q��c �E ����_t����Ë�ɋ@t��[�A��^]� �ˉA[��^]� �����������̋T$W��;t,��t��V�p�����u�+ƍH������^v3�RP���y�����_� ���V�D$Pj���!�����^� �����������V�t$��W��t�ƍP�����u�+H������v3�VP���������_^� ������̋�3ɉ�H�H�H�H�H�H�H �H$�H(�H,������������S�\$V��FW�~;�uq��    ��   v��|�  ;�}�������   ~� �V��t.��+���x%;�}!;��}Q���o���V�F���F_^[� ;�}Q����n���N��V_���F^[� �������SVW������tF��;5��t;��t7�>~2�:����FSP�������F;F}�?��t
���G_^[Ë=���G_^[���������̋D$�V��W�=����t�����3�9H����#ʅҋ�t���RPR���a���_^� �׋RPR���N���_^� ���������V�t$���W��t�������8 ~/�>$
 ��u&�����t��� ��_^� ���� ��_^� �����6;�t*��t�ƍP�����u�+H������v3�VP���������_^� ������V�������D$^� ��������������QV�t$Q���D$    �:����D$P���������^Y� �������QW�|$Q���D$    �
����T$��t��V�p�����u�+ƍH������^v3�RP��������_Y� ���V����Wt�������|$;x|W�}�����|A���t������;x,����������t���x�� _^� ����x�� _^� ���V�������6�ƅ�t��3�9H����#΋�^á��3�9H����#΋�^������̋��     �������̋��L$�� ����̋�����������������������������A�������������A������������Q��$�$�p4Y���������������Q�A�$�$�p4Y��������������Q�A�$�$�p4Y��������������VW�|$��}3�����   ~��   �t$��}3�����   ~��   �T$��}3�����   ~��   �D$��}3��=�   ~��   ���������_�^� �������S�D$U��VW��������z�����������z��������D$������z�����������Au�����D$$������z�����������Au�����D$,������z���������������Au������������x4�����������aa ���؉\$�Ta ���|$�Ga �Ë��t$$�:a �D$�ȉL$,����$��������Az���d$������u���D$$����������Az���D$,��������Az��QVWS���I���_^][�  �̋T$�ҋD$V�t$}3�����   ~��   ��}3�����   ~��   ��}3������^� =�   ~��   �����^� ���������� �\$�D$4�\$�D$,�\$�D$$�$�+���� �������̋D$�T$P�D$RP�    �F������ �U������,  ��E�M�S�VW3�h�   �T$SR��$4  Ǆ$8     Ǆ$<     ��$�   ��W ��uݔ$�   �T$t�    �T$L��$�   ��T$$݄$�   �����3�3�3ɍ�$�   �G���������Au�ً�3�������������Au�ًѾ   ����G��������Au�ًѾ   ����G��������Au�ًѾ   ��؃��� ��|��ҋE���   ��݄�   ���   ݜ$�   ���Ƀ��X���݄$�   �   �@�ݜ$�   �X�݄$�   �@�ݜ$�   �X�݄$�   � ݜ$�   ��D� ���\$���Ƀ��P��D$ �@��\$ �X��D$(�@��\$(�X��D$0� �\$0�݄$�   ����Ʌ�tn݄��   ����   ݜ$�   �� �� �X��� ݄$�   ��$(  �@���ݜ$�   �X�݄$�   �@�ݜ$�   �X�݄$  � ݜ$  �݄$�   ���$(  ����������  ݄$�   �   ��$�   ݔ$�   ݄$�   ��ݔ$�   ݄$�   ��ݔ$�   �D$���T$�D$ ���\$ �D$(���\$(�D$0���\$0������ݜ$�   ����4�T$݄$�   ����������Au��������܄$�   ݔ$�   ����܄$�   ݜ$�   ����܄$�   ݜ$�   �����D$8�T$8�D$ ���D$@�\$@�D$(���D$H�\$H�D$0�����D$P�\$P݄$�   �D$����D$8݄$�   ������݄$�   ��������Au݄$�   ������܄$�   ݜ$�   ����܄$�   ݔ$�   ����܄$   ݜ$   �������D$X�\$X�D$ ���D$`�\$`�D$(���D$h�\$h�D$0�����D$p�\$p�D$���݄$�   ��݄$  ���\$����A��   ݄$  ������܄$  ݜ$  ����܄$  ݜ$  ݄$�   ��܄$   ݔ$   �������D$x�\$x�D$ ��܄$�   ݜ$�   �D$(��܄$�   ݜ$�   �D$0����܄$�   ݜ$�   ݄$�   ���݄$   ���Ë�����\$��$�   �G����D$������z�\$�Ѿ   �������D$������z�\$�Ѿ   ����G���D$������z�\$�Ѿ   ��؃��� ��|��M��D$��������z�����   �����ڍ��   �ۃ��ۃ��ڃ�݄$�   �@�ݜ$�   �X�݄$�   �@�ݜ$�   �X�݄$�   �@�ݜ$�   �X�݄$�   � ݜ$�   ��D� ���\$8�����X���D$@�@��\$@�X��D$H�@��\$H�X��D$P� �\$P��D$8݄$   ݄$�   ݄$�   ݄$�   ݄$�   ��������������˃���   �ڍ���   �ڃ� �ڃ� �؃� �@���$,  ݜ$�   ���X�݄$�   �@�ݜ$�   �X�݄$�   �@�ݜ$�   �X�݄$  � ݜ$  �݄$   ݄$�   ݄$�   ݄$�   ݄$�   ���$,  ������������  ݄$�   �   ��$�   ݔ$�   ݄$�   ��ݜ$�   �����T$8�D$@���\$@�D$H���\$H�D$P���\$P݄$�   ����ݜ$�   �D$��4�T$����������Auj��������������ݔ$�   ݄$�   ��܄$�   ݜ$�   �����D$�\$���L$@�D$ �\$ �D$H���D$(�\$(�D$P�����D$0�\$0�D$�����݄$�   ������������Aui����������ݔ$�   ݄$�   ��܄$   ݜ$   �����D$X�T$X���L$@�D$`�\$`�D$H���D$h�\$h�D$P�����D$p�\$p݄$�   ����D$X��������݄$  ���\$����A��   ݄$  ������܄$  ݜ$  ݄$�   ������ݔ$   �����D$x�\$x���L$@܄$�   ݜ$�   �D$H��܄$�   ݜ$�   �D$P����܄$�   ݜ$�   ݄$�   ��������\$��$   �G����D$������z�\$�Ѿ   �������D$������z�\$�Ѿ   ��؃��� ��|��M��D$��������z�����   �����ۍ��   �ك��ۃ��؃�݄$�   �@�ݜ$�   �X�݄$�   �@�ݜ$�   �X�݄$�   �@�ݜ$�   �X�݄$   � ݜ$   ��D� ���\$X�����X���D$`�@��\$`�X��D$h�@��\$h�X��D$p� �\$p��D$X�D$8݄$   ݄$�   ݄$�   ݄$�   ��������˃�t~�ڍ���   �ڃ� �ك� �@��� ݜ$�   ���X�݄$�   �@�ݜ$�   �X�݄$�   �@�ݜ$�   �X�݄$  � ݜ$  �݄$   ݄$�   ݄$�   ݄$�   ���$0  �����������j  ݄$   Ǆ$�      ��ݔ$   �����T$X�D$`���\$`�D$h���\$h�D$p���\$p݄$�   ����ݜ$�   �D$��4�T$����������AuZ����������܄$�   ݜ$�   �����D$�\$�D$`���D$ �\$ ���D$h�����D$(�\$(�D$p�����D$0�\$0�D$�
���D$h��������������AuN��������܄$�   ݜ$�   ���������T$8�D$`���D$@�\$@�����D$H�\$H�D$p�����D$P�\$P���݄$  ������������AuV���������������D$x�\$x�D$`��܄$�   ݜ$�   ������܄$�   ݜ$�   �D$p����܄$�   ݜ$�   ������������������T$�����z�����������  �D$xǄ$�      ���T$x݄$�   ��ݔ$�   ݄$�   ��ݔ$�   ݄$�   ��ݔ$�   ݄$�   ����ݜ$�   �D$��4�T$݄$�   ��������AuN����݄$�   �������D$�\$�����D$ �\$ �����D$(�\$(݄$�   �����D$0�\$0�D$������݄$�   ��������AuP����݄$�   �����������T$8�����D$@�\$@�����D$H�\$H݄$�   �����D$P�\$P�D$��������݄$   ��������AuA݄$   �������������T$X�������D$`�\$`�������D$h�\$h�����D$p�\$p��������ف�  �yK���C݄$�   t���M��
���������Ƀ�t[�����D4�D4�\$X�����X����D$`�@��\$`�X��D$h�@��\$h�X��D$p� �\$p��D$8���������������	�ً�$,  ��tL���D4�D4�\$8��$(  ���X����D$@���@��\$@�X��D$H�@��\$H�X��D$P� �\$P����$(  ������؅�tG�D$���D4�D4�\$�����X����D$ �@��\$ �X��D$(�@��\$(�X��D$0� �\$0��}��$�   �    �t$�_^[��]����������������Vh�   ��j V�H ����^x��^�����Vh�   ��j V�pH �D$�����VP�V(����^x^� ������Vh�   ��j V�@H �D$�VP���V(������^x^� ������VW�|$��j ���|  �j���|  �^ j���|  �^@��|$j �^`���s|  �^j���g|  �^(j���[|  �^H��|$j �^h���F|  �^j���:|  �^0j���.|  �^P��|$j �^p���|  �^j���|  �^8j���|  �^X��_�^x��^� �̋D$��w���� 3�� ����������U������   �E� V�	W�A�H ���A�H@���A�H`���\$�@�	�@(�I���@H�I���A�Hh���\$�@�	�@0�I���@P�I���@p�I���\$�@8�I��H���A�HX���@x�I���\$ �A(�H �A ����A0�H@���@`�I8���\$(�@(�I(�@�I ���@H�I0���@h�I8���\$0�@0�I(�A �H���A0�HP���@p�I8���\$8�A �H�A(�H8���A0�HX���@x�I8���\$@�AH�H �A@����AP�H@���@`�IX���\$H�@(�IH�A@�H���@H�IP���@h�IX���\$P�@0�IH�A@�H���AP�HP���@p�IX���\$X�A@�H�AH�H8���AP�HX���@x�IX���\$`�Ah�H �A`����Ap�H@���@`�Ix���\$h�@(�Ih�A`�H�t$���@H�Ip���@h�Ix���\$p�Ah�H0�A`�H���Ap�HP���@p�Ix���\$x�A`�H�Ah�H8���Ap�HX���@x�E�Ix�    ����ݜ$�   �_^��]� ������������h�   j Q��D ������������������Vh�   ��j V��D ���Vx���VP�V(�^���������������Vh�   ��j V�D �D$����D$�^(�D$�^P���^x^� Vh�   ��j V�`D ��D$�Vx�VP���V(�� �^�@�^8�@�^X�^x^� ����U������L�E�@�Q�T$V�@ ���T$(�@(�T$0�@0�\$�@8�\$�@@�\$� �@�@3��D���L$�� �ƃ� ���L���^���L$���L���^���L$���L���^��B����B������B������\0|���^�������Q`���d$4�Y�Qh���d$<�Y8�Yp�d$D�YX���Yx��]� �������̋D$� �@�@�A��������A�����A�A(���A �����A0�����A8�AH���A@�����AP�����AX�Ah���A`�������Ap���������Ax��������D{�����������V�t$�˃��ʋ��\$�������\$���$�jr  ��^� ���̋D$� V�@�t$�@���A��������A�����A(���A �����A0�����AH���A@�������AP���������\$�\$�$��q  ��^� ���������D$3��������a���������AzZ�����������AzJ�����������Az:�����������Az*�����������Az����|��!��������Az	�� ����2�� ����3��������Dz����|��ذ���2���������������́�   ��D$P�T$�T$�\$R�D$PQ������$�   ����t�D$����$��������D{����Đ   � ���������̃�V�t$Wh�   j V���A ��D$�^x��P�L$ �\$QVW�����D$<����t�D$�_��^��� �U������   ���V�u��Q�V�A�F�Q�V�A�F�Q�V�V�A �F �Q$�V$�A(�F(�Q,�V,�A0�F0�Q4�V8�V4�A@�F@�QD�VD�AH�FH�QL�VL�AP�FP�IT�VX�V`�T$�VhR�Vp�D$��NTP�^x�L$ Q�T$V�\$�����������   �D$������4������zk����$����z^�D$������4������zI�D$��D$8�^�D$X�^�D$ �^ �D$@�^(�D$`�^0�D$(�^@�D$H�^H�D$h�^P^��]� ��������^��]� ���U������<Vh�   ��j V�g? ���Vx���VP�V(��E������4�����E��A��4z9����������Az,�������������U���������  �0'�]�  ������������u��������Az	���  ����������������������Au8�����\$�L$8�$�`{  �L$(�7q  ����   �D$(�U�D$0�U����������4�������  ������4������A�  ����������A�%���������A��������������Dz@��������Dz5����^��]�@ h�4h�4h�  h�4�eY ��^��]�@ ���U����L$(�\$�E�\$(�E �\$0�E(�\$8� s  �%�$����4����Au	�L$(�t  �D$(�����D$�����E�T$��D$0�������D$8���E�������T$ �^�������\$���T$�D$�V�������V �������E�V(�����������M�����T$(�^0�D$�d$�T$�^@�����VH�����������E�T$�^P�����E0��������D�E8z��������Dz���]@����D��   ���D$�%�$���D$ �����E@�����������^���������������D$(���������^8���D$�������D$�����������^X�������Vp�Vh�^`�^x^��]�@ �����������������������Au�0'�U���]� ������U���]�������������������������U������  VWh�   ��$�   j P����; �E� h�   ݜ$�   �L$�@j ݜ$�   Q�@�Eݜ$�   � ݜ$�   �@ݜ$�   �@�Eݜ$�   � ݜ$�   �@ݜ$�   �@ݜ$�   ��ݜ$  �r; �E� �M�U�\$ ����\$��\$�@�\$(�A�\$0�B�\$8�@��$  �\$H�A�L$�\$P�B��$�   �\$XR��Pݜ$�   ������    ���_^��]� �������U������  VWh�   ��$�   j P����: ��Eݔ$�   ݔ$�   h�   ݔ$�   ��$0  � j ��Qݜ$�   �@��ݜ$�   �@��ݜ$  ݜ$0  �t: �U$��E ݜ$�  �M��R�UP�EQ�MRPQ��$8  �4����UR�L$�j  h�   �D$$j P�&: ���T$|���T$H��$�   �T$ Q�D$��$$  �\$<R�D$��$(  �\$`P�D$$��$�  ݜ$�   Q�L$0ݜ$�   �����������    ���_^��]�  ��U�������   SVWh�   ��j V��$   �9 ��}�^x�u��V���j  ݜ$�   �]S���j  �\$S���j  �\$PW���{j  �\$X݄$�   �E�\$`P�D$���\$l�Yj  �M�\$pQ���Jj  �\$x�UR���;j  ݜ$�   ݄$�   V��ݜ$�   �j  ݜ$�   �}�D$PWݜ$�   ���j  ݜ$�   �EP����i  ݜ$�   �MQ����i  ݜ$�   �D$Sݜ$�   ���D$Tݜ$�   �i  ݜ$�   W���i  ݜ$�   �UR���i  ݜ$�   �EP���i  ݜ$�   ݄$�   �\$X����Az3���   ��    +��D�X�L$ܜ$�   ����z	�   �L$�A�   ���B�T$����4�    +�t�X�t$�����D��  ��I�����6�LX�t`�|h�\p�\$(�����������������\x����   �ɉD$,�\$$��\$���D$��D$�@���C�\�X�\�X�\$����D{m��D$���\$(��@�����DX�\X����D`�\`����Dh�\h��\$$���Dp�\p��\$,���Dx�\x���   �� ��D$����ɋ\$���R�C�\�X�\�X�\$����D{i��\$(���R������DX�\X����D`�\`����Dh�\h��\$$���Dp�\p��\$,���Dx�\x���   �� ��D$����ɋ\$��    +��D�X��    +����D�X��������Au
�Ëډ\$�Ѝ�    ��+��\�X�D�X�D$����Dz����2�_^[��]� �D$���0�[���\X�\$@�����\`��\$<����\h��\$8����\p��\$D����\x����   �ɉD$4�\$0��\$���D$��D$�@�����\�X�\�X��$�   ����D{\��D$@��� �D$<����� �D$8����� �D$D����� �D$(��� ��D$0� �D$$��� ��D$4��D$,� �����ɋ\$���R�C�\�X�\�X�\$����D{u��\$@���R��\$<�����DX�\X��\$8���D`�\`��\$D���Dh�\h��\$0���Dp�\p��\$4���Dx�\x���   �� ��D$����ɍ�    ��+��\�X�\�X�\$����D�O������R�3���\X�\$�����\`��\$L����\h��\$H����\p��\$P����\x����   �ɉD$����D$���$�   ��T�X�D�X�D$����D{\�D$� �D$��� �D$H�����L$L��L$P����� �D$(������L$��� ��D$$���� ��D$��D$,� ���D$�@�B�T�X�L�X����D{b��T$�D$@����T$H��� ��D$L� �D$<��� ��D$8��T$��� ��D$P� �D$D��� ��D$0���� ��D$4�
� ����؋�$�   �D$p�_�D$t^�X[�D$t�X݄$�   �X ݄$�   �X(݄$�   �X0݄$�   �X@݄$�   �XH݄$�   �XP���]� ������́�   ��$  ��$  VWP��$  ����$  QRP��$  �J���h�   �L$j Q�Y2 �苄$(  �T$d�T$<h�   �T$��$�   � j ��R�\$8�@���\$X�@���\$xݜ$�   �2 ��$@  �苌$<  ݜ$  ��$8  ��PQRh(�h�h����$�   � ����Ѝ�$  P��$�   Q�D$P��$�  Q��$�   �e������^�����    �_��^��   �  ��������j�h 6d�    P��SUVW�  3�P�D$$d�    ��h�   j V�D$8   2��@1 ��|$@�Vx�VP�����V(��,  j �L$<��X  �5�����D�  j�L$<��X  �5�����D��   j �L$L�X  �5�����D��   j�L$L�X  �5�����D��   �L$8�BY  ��$����D��   �D$8P�L$L��n  ����   �L$H�Y  �\$�L$8�Y  �|$j�L$<�\$ � X  j �L$L���X  � �M j�L$L�\$��W  j �L$<����W  �E ��L$8�l$�\$�X  �|$�����D$���\7�L$8�D$, 艦 �L$H�D$,�����x� �ËL$$d�    Y_^][���$ U�������  �UVW������Dz<�U����Dz2�]����Dz*h�   j W�/ �E ����W(�_P���_x_^��]�  �؍EP�L$Q��=�S`  h�   ��$�   j R���=/ ��ݔ$�   h�   ݔ$�   ��$0  ݔ$�   j �Pݜ$�   �Fݜ$�   �Fݜ$  ݜ$0  ��. �E ��ݔ$   h�=ݔ$L  �L$ݜ$t  Q��Mݜ$�  �_  h�   �T$$j R���. ���T$|���T$H��$�   �T$ P���$$  �\$<Q�F��$(  �\$`R�F��$�  ݜ$�   P�L$0ݜ$�   �����������    ���_^��]�  �����U�������|V���V`����D�   �Vh����D�  �^p����D�  ���^x����D��  j �a����T$0����4����A��  �F@���\$�L$h�F �\$��$�k]  �FH���\$�L$P�F(�\$�F�$�K]  �FP���\$��$�   �F0�\$�F�$�(]  �L$P�c  �\$�L$8�rc  �\$�L$h�ec  �T$ �����D$��������D�  ���D$��������D��   ��������D��   �������5����������   ������������A��   ������������A��   �D$8P�L$T��]  �D$�L$�L$hQ�L$<���\$,��]  �D$ �L$�T$PR�L$l���\$�]  �D$ �L$���D$(����'��������{h�D$��������AtY����������AtP���\$0����z
�   ^��]Ã��^��]���3�����^��]�����3�����^��]���3�������^��]�������3�^��]�����������̋T$(�D$V��L$(���ĉ�L$H�P�T$L�H�L$P�P�T$T�H�L$(�P�T$,���ĉ�L$H�P�T$L�H�L$P�P�T$T�H�P��? ���$�D$@�	A �����$�����^�8 �������̋D$�PHR�P0R�PRP�D$�PHR�P0R�PRP�9���� �����̋D$�PHR�P0R�PRP�D$�PHR�P0R�PRP�Y���� �����̋D$P�T!����j�h.6d�    PSUVW�  3�P�D$d�    3���9u)��9�\$��	 ����9X5t
��95�l$$�t$(3��E �E�E;�E��;���   �:�t< 
�F��:�u�>{u��3���$    3҈\$$�\$%��    ���:�td��,A<w��7�L$���*��,0<	w	�D$�����,a<w��W�L$�����-u&��|��L$$��9����L$%�����(|��#�`/�d/�h/�M �l/�U�E�M�ŋL$d�    Y_^][������������̋T$��u	�D$���ËL$��u�AËV�1;�rw#�B�qf;�rw�B�qf;�s���^�v�   ^ø   ��W�d$ �2;1u��������s��t^�2�9+�uE��������tG�2�9+�u.��������t0�2�9+�u��������t�2�+�t���   _���^�3�_^��������������������̋D$�8 u�x u�x u	�x u��2����������������̋D$�8 u�x u�x u	�x u2�ð����������������j�h^6d�    PQSUVW�  3�P�D$d�    ��9u3��9�D$     ���	 ��u�X5�5�9��5�5�9��5�9�L$,��u3��L$d�    Y_^][��Ë|$(��5��5��+�+ƍV�D$�B��48�������5������5������}� t�-���B��48�������5������5������}  t�-����4�������5������5������< t�-���B�48�������5������5����D$���< t�-���������5����� �D$,�L$d�    Y_^][�������W�|$��u
�D$���_�V�t$��u�F^_�VW���������u�G+F^_�������̋L$�ɋD$u���Å�u�   ÉD$�L$�����������̋D$��v	�D$�E6 3�������������̋L$��v�D$��v�D$�L$�KI 3�ËD$��t	�D$��6 ��������������̋D$��w�D$��t	P�6 ��3�ËL$��u
P��5 ��ÉD$�L$�,I �����V�t$��th�9��������t��^�3�^���������������̸�9�����������Q�`/V��F�d/�N�h/�V�l/�F�`/�N�d/�V �h/�F$�l/W����N(�N4�~�~,�~0�� j j j �NH�~D������`/�VL�d/�FP�h/�NT�l/W�L$�VX�$�����D$�^`�Nh�F\�P� �_�Fl�Fm �Fn�Fo ^Y������������̃�h�H� ��t�D$��th�5P��� ��3�� �   � ̸@   ����������̋D$V��P�Nh�� ��Bj ���Ѕ���^� �����������̋D$V��P�Nh��� ��Bj ���Ѕ���^� �����������̍Ah������������̋D$�AH� �����̋IH�D$�� ���̊Al������������̊Am������������̀yl t�ym u�   �3������������̋A0�������������VW��V3���������uy�N��������t�   �N�������t�����^����A{�F�0'����Dz�F���$�J  ����t���F <t<u���F!<t<u�� ��t����_^����������������Q3�V���F�F�F�F�F�F�F�F j��L$�F$�����D$j��L$�F������5�L$�^�N^Y��������������VW�|$jj��h � @���h� ��u_^� S��2�������D$�D$Pj���� ����   �|$ ��   V���� ����   �D$   t�NQ���;� ��t}�D$   t�VR���"� ��td�D$   t�F�����$��� ��tF�D$   t �F P���
� ��t,�N Q����� ��t�D$    t�V!R����� ��t����� ��u2ۊ�[_^� ����̃�UVW�������|$�D$P�L$Q3�h � @�ωl$�l$�/ ��u	_^]��� S2ۃ|$��   �T$ Rj�ωl$(�� ����   9l$ ��   V���� ����   �   �l$ t�FP����� ����   �D$    t�NQ����� ����   �D$    t�VR���� ��th�D$    t%�F P���G� ��tO�|$|�N!Q���1� ��t99l$|�D$     t�V!R���� ��t�D$��P��������t�F! ����-
 ��u2ۊ�[_^]��� ����������̸�:����������̋L$h 6�� �   � �����������˱�������������V��踱���D$t	V�K�������^� ��QV��j �L$ǆ�       ������D$j �L$���   �������L$ݞ�   ���   Ɔ�    Ɔ�    ^Y���������������̸�;�����������VW�|$W���w ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ݇�   _ݞ�   ��^� ���j�h�6d�    P��V�  3�P�D$d�    ��t$�Av ���   �D$$    �d6��������   ������D$P��;�^�����N�P�V�H�N�P�V� 0�F�0�N�0�V �0�ΉF$�F(   �����ƋL$d�    Y^�� ����̸   � �������̸�   ����������̋D$VW�񍾸   WjP�6 ������t���   RjP��5 �������t���   RjP��5 �������t���   RjP��5 �������t���   RjP�5 �������t���   VjP�5 ��_^� ������VW�|$j j��h � @���8{ ��u_3�^� ���   SP��2��� ����   ���   ����t���   R���)� ����   ���   ���t���   Q���� ��th���   ����t���   P���u ��tG���   ����t���   R���T ��t&���   ���t݆�   �����$�� ��t����� ��u2���[_^� ���̃�UV�������l$3��D$�D$�D$P�L$Qh � @��� ��u
^3�]��� S2ۃ|$��   W���   W���u� ����   �����t���   P����� ��tq�����t���   R����� ��tU����t���   Q���� ��t:�����t���   P���c� ��t�����t���   V���w� ��t�_���Y ��u2���[^]��� ������̋��   ��>�����ËL$h�6��� �   � ����������V��FP�t�������t�|$ �No������   
ȈNo^� �No2����
ȈNo^� ��������������VW�|$��;~teS3�;�~D9~~�~�N��PWQ����;ÉFt:�N;�~��+���R���SQ�D ��[�~_^� �F;�t�SP�B�Љ^�^�^[_^� ��������̋A��~�I���D���3�������������j�h�6d�    PQ�  3�P�D$d�    �L$�L$���D$    t�6� �L$d�    Y��� ����VW�|$��;~tlS3�;�~K9~~�~�N��PWQ����;ÉFtA�V;�~��+ʍ����Q����SP�M ��[�~_^� �F;�t�SP�B�Љ^�^�^[_^� ��SW�|$����~dU�l$��|ZV�t$��|P;�tL�C�/;�B;�>�K�>;�~�;�}��P���6����C�����R�L� ��R����R�5 ��^]_[� �����������SVW���Oh�� �؅�u��7�G�t$Ph�7V��� Sht7V��� ���l �l7u�d7PhT7V�� ���m �L7u�@7Ph07V�� h7V�� ���OHQ���� h�&V�w� h7V�l� ���W\R���� h�&V�S� �G0Ph�6V�D� ��_^[� �����������QV�t$Wj��j���� ����  �l Su)�GP�4�������t�Go����t	��u2�����_l�m �\$t)�OQ���������t�Go����t	��u2�����Gm�ۈD$[t3��3҄�����P����� ���\  �GP���� ���I  �O,Q���� ���6  �W0R���� ���#  j ���� ���  �GHP���� ����   j ���� ����   j ���� ����   ������$��� ����   ������$�� ����   �OhQ���� ����   �T$R���6� ����   �GDP����� ��ty�O\Q���� ��tj�G`�����$�`� ��tV�T$R����� ��tF�GP���� ��t7�OQ���� ��t(�WnR����� ��tV�O4�%� ��t��LW���V� _��^Y� ������������̃�S3�UW���\$�\$�\$�\$�A����l$(�D$P�L$Q����� ��;���  �|$�x  V�T$R����� ��;��;  �D$+Í_lt��t���u�Gm�� ���Gm �GP���� ������  �O,Q���� ������  �W0R���� ������  �D$P���v� ������  �OHQ��� � ������  �T$,R��詿 �D$,P��蝿 �L$ Q����� �T$ R���� �GhP���
� �����\  �|$�Q  S���\� �����>  �|$�3  �ODQ���ۿ �����  �|$�  �W\R���Z� ������   �G`P���4� ������   �|$��   �GmP����� ������   �|$��   �OQ���� ������   �|$|m���	-	 =w�~_�GP���W� ����t}�wV��������t/�; tV�����Wo����������
ЈWo�m u	j ���a����GnP���F� ����t,�|$|%U�O4�� ����t�|$|�OLQ����� ����W�j�������t	W���������^_][��� h�7h�7h�  h�7�%. ��_]3�[��� �������S�\$V��W�����~W�Fl��������t
�fo�_^[� ��tW�����No����������
ȈNo_^[� S�\$V��W�����~W�Fm��������t
�fo�_^[� ��uW������No���������
ȈNo_^[� S�\$VW�|$WS�^�����������   U�������ϋ�������+���   ��   t�s �G +���   ��    t�s!�O!+�um��   t�K�*����O��� ���+�uO��   t�K�����O������+�u1��   t)�G�[����Au
]���_��^[��G�[����z�   ]_��^[�������VW�|$��tMh�:���ʝ����t=�t$��t5h�:��貝����t%W���i ���   �P���   �Ǹ   W��_�^�_2�^����̋��   ����   ���������������̋��   ���   ����P�Qj ��( ��� �����������̃�SVW�|$j ��jh � @�ωt$�n �؄�u_^3�[��� ����k ���D$t`h�9��������tPU���   U����� �؄�t:3���~43��I ��t'�D$���   �T$�D$R�P��������(;���|Ջ|$]���y� ��u2�_^��[��� �������SU�鋝�   V3���W~)3��
��$    �I ���   ��C�����u����(;�|�_^]�[�_^]2�[��������j�h�6d�    PQ�  3�P�D$d�    h�   �������D$���D$    t���{����L$d�    Y���3��L$d�    Y������������j�h7d�    PQVW�  3�P�D$d�    ��h�   �������D$���D$    t���������3����D$����tW�������ƋL$d�    Y_^������������VW�|$��t5h�;��������t%�t$��th�;��������tW���6���_�^�_2�^�������������V���d6�"g �D$t	V���������^� ������������S�\$��VW��}%�F3�;���   �WP�B�Љ~�~�~_^[� �F;�}v��F�RSP��3�;ǉF�   �VU��+ʋ���+������U+ʍ�WR� �F��;�}$����+�����+�F�P���r�����<��u�]_�^^[� ~&9^~�^��F�RSP�^��3�;ǉFu�~�~_^[� ��V��~ ��6t%�F��tj P��6�F    �F    �F    ^�����������V��L$��|H�F;�}A+���P�APQ�������F��N�V3����ʉ�A�A�A�A�A�A�A�A �A$^� ���������V��~ ��6t%�F��tj P��6�F    �F    �F    �D$t	V���������^� ������j�hV7d�    P��V�  3�P�D$d�    ��t$��c 3��8�D$$ǆ�   �6���   ���   ���   �D$P��:�D$(�Օ����N�P�V�H�N�P�V� 0�F�0�N�0�V �0�F$�F(   �ƋL$d�    Y^�� ���j�h�7d�    PQSVW�  3�P�D$d�    ���|$�83�9��   ���   �\$��6t�F;�tSP����6�^�^�^���D$������c �L$d�    Y_^[��������������������������V��FW3�;��H8tWP�T8�~�~�~_^���������̋Q2���t%�I��~V�t$��t��~Vj<QR�{ ���^� ��������������̋Q2���t%�I��~V�t$��t��~Vj<QR�h{ ���^� ��������������̋D$�T$����+���QR�F������ ���  3ĉD$SV��F�V;�W�|$$��   ������   v��|� � ;�}�������   ���^��tD��+���x;;�}7;ЋO�U�o��L$}P��������F�T$��F��h�P�x]�+;�}P��������F���F��W�P�O�H�W�P�F�L$_^[3��~ ��� ��������������SU�l$��;�tT�E��]�C    ��[� 9C}P������{ t.�E3҅��C~"V3�W�u�{���   ����<;S|�_^]��[� ���������V��F���H8tj P�T8�F    �D$�F    �F    t	V�%�������^� ������������V��F�V;�u?����Ɂ�   v��|�;33 ;�}�������   ��;�}P���d����N3����N�щ�A�A�A�A�A�A�A�A �A$�N�F�����N��^������j�h�7d�    PQSVW�  3�P�D$d�    ���|$�\8�wh���D$   �>� ���D$�2� �G8�w43�;È\$�H8tSP���T8�^�ω^�^�D$�����Z����L$d�    Y_^[����������j�h�7d�    PQ�  3�P�D$d�    h�   �������D$���D$    t�������L$d�    Y���3��L$d�    Y������������j�h+8d�    PQVW�  3�P�D$d�    ��h�   �A������D$���D$    t���7������3����D$����t W����^ ���   �P���   �Ǹ   W�ҋƋL$d�    Y_^����j�h[8d�    P��VW�  3�P�D$ d�    �D$P��:������|$0P��耐������th�:���~�����uB3�8D$8tUh�   �x������D$���D$(    t���n������3�V���D$,����踗���D$4� ��ƋL$ d�    Y_^�� ËL$4�	�L$ d�    Y_^�� �����V��������D$t	V���������^� �̃�SUVW�����   3�9^|�^�l$ �D$P�L$Qh � @�͉\$ �\$$�� ��u_^]3�[��� ���n` ��;�th�9���|�����u3�;��Ä���   �|$�Ä���   �T$R���D$    �E� �؄���   �D$9F}P��������D$3��~W�D$ PW�������������؄�t-���?������������u�F��R��P���҃�;l$|���N��P��Q����h�~����J �l$ ���2� ��u2�_^]��[��� ��������������̃� �  3ĉD$�L$0�D$,�T$4SUV�t$0�L$W�|$8�D$�D$H�L$Q�T$(�D$,���������)  �T$LRWV�e���������  ���   ���   3����D$�L$��   �L$��    �   �T$��$    �2;1u��������s��t]�2�+�uE��������tF�2�+�u.��������t/�2�+�u��������t�2�+�t���   ����3����&  �L$����(;|$�L$�Y����|$L �6  ���   ���A������   ���Ήl$������D$��L$ �N�T$$�V�D$(�F�G��t&���~��~��t��~h�~j(WP�is ��3�9\$��   �����    �   �ύT$��I �2;1u��������s��tz�2�)+�uE��������tc�2�)+�u.��������tL�2�)+�u��������t5�2�+�t+���   $�����T$��_^]��[�L$3���� �� �3���t%����(;\$�H���_^]3�[�L$3��� �� ËL$_^�����L$$][3��� �� �������VW�|$W��袘���G�F�O�N�W�V�G�F�O�N�W�V�G �F �O$�N$�W(�V(�G,�F,�O0�W4�N0R�N4������GD�FD�OH�NH�WL�VL�GP�FP�OT�NT�WX�VX�G\�Oh�F\�G`Q�^`�Nh��� �Wl�Vl�Gm�Fm�On�Nn�Wo_�Vo��^� �������VW�|$��t5h�9���
�����t%�t$��th�9��������tW������_�^�_2�^�������������j�h�8d�    PQV�  3�P�D$d�    ��t$�C����N4�D$    �\8�]� �NH�D$�@����N\�8����Nh�`� ���D$�Fo �p����ƋL$d�    Y^����������������V��������D$t	V�;�������^� �̃��D$�PSUV���L$�H�T$�P�D$WP�L$�T$ ��������j tX�NoQV����������}   ���   3���~q3����   �������u����(;�|�2�_^][��� �_^][��� �T$�L$���ĉ�T$,�H�L$0�P�VoRV�H���������t���U�����u�_^]2�[��� �����j�h�8d�    PQ�  3�P�D$d�    jp�(������D$���D$    t���.����L$d�    Y���3��L$d�    Y���������������j�h�8d�    PQVW�  3�P�D$d�    ��jp贽�����D$���D$    t���������3����D$����tW�������ƋL$d�    Y_^���������������V�t$��th�<���;�����t��^�3�^���������������̸�<����������̃�SV�t$W���D$P�L$Q���D$    �D$    �ÿ �؄�t	�|$t2ۄ��D$���  �WR���ܪ �؄���  �G P��觨 �؄���  �L$Q���Ѧ �؄��x  �D$���l  <u7�WR���\� �؄��S  �D$P��薦 �؄��=  �D$���1  <u7�OQ���!� �؄��  �T$R���[� �؄��  �D$����  <u7�G$P����� �؄���  �L$Q��� � �؄���  �D$����  <u7�W(R��軧 �؄���  �D$P���� �؄���  �D$����  <u5V�O,�� �؄��i  �L$Q��謥 �؄��S  �D$���G  <u7�WPR���� �؄��.  �D$P���q� �؄��  �D$���  <u7�OTQ��謧 �؄���  �T$R���6� �؄���  �D$����  <u7�G`P���a� �؄���  �L$Q����� �؄���  �D$����  <	uI�T$R���դ �؄��|  �D$P��� ���L$Q�ΉGh认 �؄��U  �D$���I  <
u7�WlR���I� �؄��0  �D$P���s� �؄��  �D$���  <u:���   Q���k� �؄���  �T$R���5� �؄���  �D$����  <u:���   P���� �؄���  �L$Q����� �؄���  �D$����  <u:���   R���ϣ �؄��v  �D$P��蹣 �؄��`  �D$���T  <u:���   Q��董 �؄��8  �T$R���{� �؄��"  �D$���  <u:���   P���S� �؄���  �L$Q���=� �؄���  �D$����  <u:���   R���� �؄���  �D$P����� �؄���  �D$����  <u:���   Q���ע �؄��~  �T$R����� �؄��h  �D$���\  <u:���   P���� �؄��@  �L$Q��胢 �؄��*  �D$���  <uL�T$R���]� �؄��  �D$P�� ���L$Q�Ή��   �3� �؄���   �D$����   <u7�WpR���� �؄���   �D$P����� �؄���   �D$����   <u.���   Q���� �؄�t{�T$R��辡 �؄�ti�D$��ta�|$ ~:<u+��XW���Z� �؄�tE�D$P��舡 �؄�t3�D$��t+�|$~<w ��th�9h�9h�  hp9�� ��_^��[��� ����W���GP��������t�D$��th$:P蚵 ��3�_� V�t$V�O,�� ��u��th�9V�p� ��^3�_� ^�   _� ���������������   %  �yH���@P�'� ���������   %  �yH���@P�� 3Ƀ����������������̊��   �������������   ��P�Ь ������������������   P賬 ���������������������   P�� �����������������̋D$VP���� �����   ^� ������VW�|$��;~tkS3�;�~J9~~�~�N��PWQ����;ÉFt@�N;�~��+�iɘ   iҘ   R�SQ�� ��[�~_^� �F;�t�SP�B�Љ^�^�^[_^� ���V��F��t�N��Qj P�g� ���F    ^������������VW�|$��;~teS3�;�~D9~~�~�N��PWQ����;ÉFt:�N;�~��+���R���SQ�� ��[�~_^� �F;�t�SP�B�Љ^�^�^[_^� ���������S�\$��U��~[W�|$��|QV�t$��|G;�tC�E�;�9;�5�M�;�~�;�}��P���6����E����S����WV��� ��^_][� ����j�h19d�    PQ�  3�P�D$d�    �L$�L$���D$    t�� �L$d�    Y��� ����SV�t$W�   S��j���h� ���E  �GP��腲 ���2  �O Q��肰 ���  U�o��蟯 ��u S���3� ����  U���� ����  �o���q� ��u!j���� ����  U���Գ ����  ���9o$t$j���ۭ ����  �W$R����� ����  9o(t$j��貭 ���~  �G(P���ϯ ���k  �D �4 8_Lu8_Mu�O,�I� ��t"j���l� ���8  V�O,苀 ���'  �oP���Y�����t!j���<� ���  U���� ����  �oT���*�����t!j���� ����  U���ݰ ����  �G`��$����D{)j���ܬ ����  �G`�����$蔰 ����  �h t,j	��譬 ���y  �Oh�L$�T$R��蒬 ���^  9_lt$j
���|� ���H  �GlP��虮 ���5  8��   t(j���P� ���  ���   Q���� ���  ���    t(j���� ����  ���   R���� ����  ���    t(j���� ����  ���   P���׫ ����  ���    t(j��轫 ����  ���   Q��覫 ���r  ���    t(j��茫 ���X  ���   R���u� ���A  ���    t(j���[� ���'  ���   P���D� ���  ���    t(j���*� ����   ���   Q���� ����   ���    ~'j����� ����   ���   R���s� ����   9��   t+j���ʪ ����   ���   �D$�L$Q��謪 ��t|�_pS��������uj��菪 ��t_S��裮 ��tS���    ~j���m� ��t=���   R����� ��t+�X tj���H� ��t�GXP���i� ��t	j ���,� ]_^[� �����QV�t$W�����u ��|V���s���_��^Y� jj���߱ ����  �GP����� ����  �O Q����� ����  �W(R���� ����  �GPP��胭 ����  �GhP���� ����  j ���� ���|  ������$�7� ���e  ������$� � ���N  �OlQ���m� ���;  ���   R���&� ���$  ���   P���� ���  ���   Q����� ����  ���   R���� ����  �GP��议 ����  �OQ��蛮 ����  ���   R���5� ����  ���   P����� ����  ���   Q���� ���v  �WhR��蕪 ���c  ���   P���N� ���L  �OTQ���� ���9  ���   R���$� ���"  �G`�����$�ܫ ���
  �G$P���)� ����   ���   �� �D$ t��t��u�D$��D$ �L$Q��迧 ����   U���   ��l$}�D$    �l$���   Su�WpR�y�������u��E�2ۋ�P��蟩 ��t��t�GpP���|� ��thP9���l� 3�;�\$~9����t@���   �U���L� ��t��U���=� �L$���� ;L$�L$|Ʉ�t	V�O,�,z []_��^Y� �SVW�񋾘   ��N��	� �N����� ؋΍��   ��y����_^[�������̋D$SVP��肢 ���   ��Q���p� ����Ã����   ���   ^[� ̀|$ V����8��   t:���   ���   %  �yH���@P�� ����t3�8��   ��Q���s���^� ���������������V�t$��P���   Q���ҋF^� ����V���   3�3҅�~*���   W�|$��    99t����;�|�_^� �   _^� ��̋��   ��~���   �D����t� Ã����V��~ �d:t%�F��tj P�p:�F    �F    �F    ^�����������S�\$��U��~dW�|$��|ZV�t$��|P;�tL�E�;�B;�>�M�;�~�;�}��P�������Eiۘ   i��   i��   S��WV��� ��^_][� �����������VW�|$��;�tA�G��_�F    ��^� 9F}P�$����N��t�G�Fi��   P�GPQ�� ��_��^� ������������V��L$��|9�F;�}2+���P�APQ��������F��Fi��   Fh�   j P�� ��^� ��������V��~ �P:t%�F��tj P�\:�F    �F    �F    ^�����������V��L$��|?�F;�}8+���P�APQ���l����F��N3���N��A�A�A�A�A�A�A^� ��V��F�V;�u;������   v��|� @ ;�}�������   ��;�}P���x����F3���F��H�H�H�H�H�H�H�N����F���N^����V��~ �d:t%�F��tj P�p:�F    �F    �F    �D$t	V��������^� ������V��~ �P:t%�F��tj P�\:�F    �F    �F    �D$t	V迩������^� ������QSVW���Er���`/�F�d/�N�h/�V�l/�N�F�{� �N�s� ���3ۍN,�^ �F$�F(�}� SSS�L$�!����SS�NPS�L$�������^`���   �VT�^X�^h�Fl   ���   Ɔ�   ���   ���   ���   ���   ���   9_t�G;�t�SP�B���Љ_�_�_ǆ�      �`/�Np�d/�Vt�h/�Fx�l/�N|�Ɯ   9^t�F;�t�SP�B���Љ^�^�^_^[YÃ�VW��������t$$���l ��|!��� 	 =���|V���.���_��^��� SU�D$P�L$3�Q�Ήl$ �l$��� ���\  �|$�Q  �WR���� �؄��  �G P���� �؄��j  �O(Q���Α �؄��U  �WPR���Y� �؄��@  �D$,P�Ήl$0��� �؄��&  ����k ��|���B� =�o�}�L$,��Q讝 ���Gh�T$,R��輐 �؄���   �D$ P���֑ �؄���   �L$ Q����� �؄���   �WlR���� �؄���   ���   P���C� �؄���   ���   U���+� �؄�tv�M Q苛 �E �����   U���� �؄�tR�U R�כ �E �����   U���� �؄�t.�E P賛 ���OQ�ΈE �r� �؄�t�WR���a� �����   %  ����   yH���@P� � �������ۈM ��  �|$��  ���   R��賗 �؄��i  �|$�^  U���f� �؄��L  �|$�A  ���   P���C� �؄��)  �|$�  �D$P���D$     躏 �؄��   �L$Q�� �����   U�ΉGh�ҍ �؄���  �U R�.� �E ���GTP���� �؄���  ���   U��蕍 �؄���  �M Q�1� ���W`R�ΈE ��� �؄��v  �|$�k  �G$P���� �؄��V  �|$�K  �L$,Q���D$0 �*� �؄��0  �T$,���ڍ��   ��҃����   �����D$P���D$    諎 �؄���   �D$����   P�������|$ �D$     ��   ����   ���   ������U���}� �؄�tY�EP���l� �؄�tH�EPhP9��������u3�M �Op�U�Wt�E�Gx�M�O|���   ���   �R���   ��P�ҋD$ ��;D$�D$ �o������    u���   �5! ��t!�|$|V�O,�1� ��]��[_^��� 2�]��[_^��� ���SUVW���O�� ��u��7�t$Ph4;V�9� h$;V�.� ���GP��耦 h�&V�� ���   ��  �yI���AQ�� ���� t��t��t�,1��L7��d7��;Ph;V�ß �W Rh�:V负 �G(Ph�:V襟 ���   Q�,1�� ��(�� t��t��u��:���:���:Sh�:V�b� ���   ����~O���   h|:V�D� ��3ۅ�~'��t��Rhx:��Pht:V�� ����;�|�h�&V�	� ��_^][� ��������������̋D$��V��|P�������u�D$P���   苁��^� ������̃��    V���   t(�F��t!�j P�B�����F    �F    �F    ^�������S�\$��UVW��}o3�9~t[�^��xB�����F�|( �|(�d:t�G��tj P���p:3��G�G�G���� ��}�3���F�RWP���҉~�~�~_^][� �F;�}m�N��PSQ����3�;FtI�N��+���W��R�Q�]� �F��;�}������+�F�P��������� ��u�_�^^][� _�V�V^][� ~���;�|P��+������D$��$    �N�|) �|)�d:t�G��tj P���p:3��G�G�G�� �l$u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� ������j �P;�s�����̋Q2���t%�I��~V�t$��t��~Vj QR�O ���^� ���������������U�l$V��;�ty�ES3�;��^[��^]� 9F}P����9^t�E;ÉF~�W3����E�N�8ǉ9�PωQ�P�Q�P�Q�Q����P�B�Ѓ��� ;^|�_[��^]� ��^]� ����V��j �P;�����D$t	V�S�������^� ����������j�hX9d�    PQVW�  3�P�D$d�    ��t$3��NW�|$�P;�2����F;��D$�����H8tWP���T8�~�~�~�L$d�    Y_^�����������j�h�9d�    PQSVW�  3�P�D$d�    ���|$�d;���   3�9^�D$   �P:t�F;�tSP���\:�^�^�^9��   ���   �D$��$t�F;�tSP����$�^�^�^�O,�D$������O�D$�� �O�\$�� ���D$�����Sn���L$d�    Y_^[���SUVW�|$W���s���G�F�O�N�W�V�G�OQ�N�F�L� �WR�N�@� �G �F �O$�N$�W(�_,�n,S�͉V(�����CP�M�t����K �M �S!�U!�C"�E"�K#�M#�WP�VP�GT�FT�OX�NX�G`�^`�Wh�Vh�Gl�Fl�Op�Np�Wt�Vt�Gx�Fx�O|�N|���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   �R���   ���   ���   ���   ���   P�ҋ��   �P���   �ǜ   W��_��^][� ���������������VW�|$��t5h�<���:g����t%�t$��th�<���"g����tW���F���_�^�_2�^�������������j�h%:d�    PQVW�  3�P�D$d�    ��t$�rd��3��N�|$�d;讕 �N�D$衕 �N,�D$�4� �NP�D$�W~���NT�O~��ǆ�   �$���   ���   ���   ǆ�   P:���   ���   ���   ���D$�����ƋL$d�    Y_^����������V���x����D$t	V�+�������^� ��j�hK:d�    PQ�  3�P�D$d�    h�   ��������D$���D$    t��������L$d�    Y���3��L$d�    Y������������j�h{:d�    PQVW�  3�P�D$d�    ��h�   聘�����D$���D$    t���W������3����D$����tW���m����ƋL$d�    Y_^�������������5�\$����D{�D$
%�  f=�t�   �3����������5���P����3�9D$����� �3�9D$����� ��5���D$��������D{!�D$
%�  f=�t�������	�A����� ��� ����5���D$��������D{E�D$
%�  f=�t6����A�����D{!���A������Dz����� �!�A�!��� ��� ��� ����������������5�����D{.f�Af%�f=�t �Y����D{f�Qf���f���t�A�!���������������������A�����Au<�5�����D{+f�Af%�f=�t�Y����D{f�If���f���t����2��������A�����z<�5�����D{+f�Af%�f=�t�Y����D{f�If���f���t����2��������A�����D{<�5�����D{+f�Af%�f=�t�Y����D{f�If���f���t����2��������5�����D{.f�Af%�f=�t �Y����D{f�If���f���t�   ���3�����������������52����D$��������D��   �D$
%�  f=���   �������D��   f�Af%�f=�t{���Y����D{qf�Af%�f=�tc�A�����u3���   �|$ ��    �
��t!��Au+��Y����z	���� ��2Ҋ�� ��u�+��Y����Az���� ���؊�� ���������������VW�|$�j ���$���	�����tQ�Gj �����$�������t;�|$ S�t8�j�����$�������u#�Gj�����$������u[_^� _2�^� ��[_^� ������5�����Dz�Y����D{����A����Y�������A����Y����������A��Y�����̋T$�BV��W��������B����z?��������Au�ٸ   ��3��B�a�����B��A�   z
�B�p3��N�3��~�E��������Au�ظ   ��3��B�x���%�������Au�B3��p�x�3��x�B�   ������������_^����D{�� 2�� ������������̋T$��tI�B`�	�Bh�I���Bx��������D{�����B �	�B(�I���B8���B�I��	���B������Y� �����������̋T$��t~�B`�	�Bh�I���Bp�I���Bx��������D{�����B �	�B(�I���B0�I���B8���B@�	�BH�I���BP�I���BX���B�I��	���B�I���B������Y�Y� ��������D$����D$�X� �������������̃|$ ��~��� ̋��L$���A�X�A�X� ������̋��L$��~��|��� ��� ������D$����D$�X�D$�X� ������̋��L$��t���A�X�A�X� ���P�P�� �����̋��L$�� ��A�@�X�A�@�X� ��������������̋D$����\$�D$� ��|�A�\$�D$� �A�\$�D$� �������������Q�Q������������A���Y�A���Y���������̋��������������̋��L$��t���A�X� ���P�� ��������������̋��L$���A�X� ������������̋��L$�� ��A�@�X� �������̋T$������Dz�B�Y����Dz2�� �� ���������̃|$ ��~��� ��D$����D$�X�D$�X� ������̋��L$���A�X�A�X� ������̋��L$���A�X�A�X� ������̋�� �D$������@���X�H�X� ̋��L$�� ��A�@�X�A�@�X� ��������������̋��L$� �!��@�a�X�@�a�X� �����������������D$�D$������A���X�I�X� ��������������̋T$��D$���B�A�X�B�A�X� ������������̋T$��"�D$��A�b�X�A�b�X� ������������̋D$�@�I� �	���@�I��� ����̋T$������Dz�B�Y����Dz�B�Y����Dz2�� �� ����������������Q�Q������̋L$��D$�D$������A���X�I�X�������������̋��L$���A�X�A�X���X� ���D$���T$�D$��������Au�T$����;������z������$�� �L$�����������z�D$
%�  f=�t�������������������A���\$��$�|�������������������A���Y��U������<V���F���\$��$�@����T$0���D$&��%�  f=���   ��;������z�ذ�����~�^^��]���������z{�؃����;�����T$@�F�����T$H�\$�$������T$0���L$&���  f���t%��;������z�D$0�����|$8�^^��]���2�����^^��]����2��^^��]����������������������Dz�Y����Dz�   ���3�Ë��L$��t���A�X�A�X� ���P�P�� �����̋��L$���A�X���X� ����������D$����A���X�A���X� �����D$�t$�����A���X�I�X� ��������������̋T$������Dz�B�Y����Dz�B�Y����Dz�� 2�� ������������̋D$���� ��|�A� �A� �̋��L$��~��|��� ��� ������A�����������z���A��������At�   ����A��������Au�   �3���������������������A��������Au������A��������Au�����������A��A�������������������������D$���T$�D$���D$����������u������u�T$���������uB������u9�T$��������;������z&������������$��������� �L$�������������������z�D$
%�  f=�t����������������A���\$�A�\$��$�5������������A���Y�A���Y����������U������<V���F���\$�F�\$��$������T$0���D$��%�  f=���   ��;������z�ذ�����F���^�~�^^��]�����������   �؃����;�����T$@�F���T$H�F�����T$P�\$���\$�$�W����T$0���L$���  f���t.��;������z�D$(�����D$0���^�|$8�^^��]���2�����V�^^��]����2��V�^^��]������������������D$��������u$�A��������Az�A��������Az
�   � ��3�� ���������Dz�Q����Dz�Y����Dz�   ���3���������5�����D{M�Q����D{C�Y����D{;�A���\$�A�\$��$�2����%�$������4����Az�   ���3����������������̋D$�L$�@�I� �	���@�I�����̋T$�L$�B�I�D$�A�J����A�
�B�	���X�B�	��I���X�������5�����D{Cf�Af%�f=�t5�Q����D{+f�Qf���f���t�Y����D{f�Af%�f=�t����2������������5�����D{+f�Af%�f=�t�Y����D{f�If���f���t����2�����5��������Dz�A������Dz�A������Dz�   ���3�������������D$��D$�Y� �D$��D$�Y�D$�Y� ����������D$��D$�Y� �D$��D$�Y�D$�Y� ���������SV��L$2�������tw�L$$������tj�D$$����D$D�V�D$L�V�\$�\$�$�������������;����Au	����������F�L$��L$���F�L$�����^^[�0 ^��[�0 ��������������������P�P�X��5�����D{`f�Af%�f=�tR�Q����D{Hf�Qf���f���t8�Q����D{.f�Af%�f=�t �Y����D{f�If���f���t�   ���3���������������A�L$��L$���A�L$���A� ���A�������   �5�����D��   f�Af%�f=���   �Q����D��   f�Qf���f�����   �A �Y����uw�Q����D{mf�Af%�f=�t_�Q ����D{Uf�Q&f���f���tE�A(�Y����u8�Q����D{.f�Af%�f=�t �Y(����D{f�I.f���f���t�   ���3��VW�|$h,<W���� ����������uh <W�� ���F(��0�\$(�F�\$ �F �\$�F�\$�F�\$��$h�;W�ˁ ��8_^� ����D$����D$�X� ���������������A�����zF�5�����D{5f�Af%�f=�t'�Y����D{f�Qf���f���t3Ұ���������3�2����������5��Y������A�����zF�5�����D{5f�Af%�f=�t'�Y����D{f�Qf���f���t3Ұ���������3�2����������A�����zF�5�����D{5f�Af%�f=�t'�Y����D{f�Qf���f���t���A��Y����������������̋T$������Au�������� ������z�   ����� �B�Y����At��B�Y����{�3������ ���������̋T$������Au�������� ������z�   ����� �B�Y����At��B�Y����{�3������ �����������5��SV���2�W�|$ ����Dz�V����Dz�����Dz
�W����D{u����������\$������D$������u����؋��\$�����\$�������D$������Az������D$������Az�_��^^[��� �����5�_�^^��[��� ��5��S��U�l$ VW�|$$�2ۋ�����Dz�W����Dz�U ����Dz
�U����D{x���������\$��������D$������u����؋��\$�L����\$���A����D$������Az������D$������Az�_��^^][��� �����5_��^^]��[��� �����U������4SV���FW�}���\$3��F�\$��$������\$P�G�\$�G�\$��$������L$P����������zc���F�O���G�N�����\$8�E�� �D$8������u�ٍC��_^[��]� ����������u���_^[��]� ��_^[��]� _��^��[��]� ����U������tS�]VW����������   �}����������   �u���v�����t~�C���\$�C�\$��$������\$P�G�\$�G�\$��$������\$X�F�\$�F�\$��$������4���D$8������A{�D$@������Az��������2�_^[��]���������Az��2�������_^[��]����������T$8�������T$@�����T$H���G�K���C�O�������G�N�����F�O�����������C�N���C�N������������������At+����������At������������At�����ذ_^[��]����`<��������A������������������������������W�D$TSP�����D$L�L$D��P���L$t�$Q����� �@���@������N���N���L$H���%�$����4����A�����V�T$lWR�H����D$T�L$L��P���D$\�$P�<���� �@���@�C����������K���L$8���%�$����4����A�<���S�L$lVQ������D$T�L$D��P���T$\�$R������ �@���@�G����������O���L$@���%�$����4����A�����_^2�[��]����S�\$V�t$W�|$SWV���������u_^2�[��F���\$�F�\$��$�!����%�$������4����At��G���\$�G�\$��$������%�$������4����At��C���\$�C�\$��$�����%�$������4����A�]���_^�[����������S�\$V�t$W�|$SVW��������u_^2�[��G�N�F�O����O��N���F��G����C����������K����4����A{�_^�[�̋D$��A�A�@ ��� �����@@�����@`�@(���@�����@H�����@h�@0���@�����@P�����@p�@8���@�������@X���������@x��������D{���������D$��������������X���X� ����̋T$��"�D$��A�b�X�A�b�X� �������������SV���F���\$2��F�\$��$�/������������z������F���^�~�^^[�^�؊�[�̋T$��"�D$��A�b�X� �����̋D$�@���a�\$�@�a�\$� �!�$������� ���U������   ��E�UV���V�M�V�� �!�\$0�@�a�\$8�@�a�\$@�� �T$�B�`�T$ �B�`�T$(��"�T$H�A�b�T$P�A��$�   �b�T$X������������������������������ݜ$�   ݜ$�   ݜ$�   �������u	2�^��]� �D$P�L$`���D$@���D$X���D$8�������D$0���D$H�������������������\$`���\$h�\$p������t��D$(��$�   ���D$8���D$ ���D$@�������D$���D$0����������������ݜ$�   ��ݜ$�   ݜ$�   �2������C����D$@���\$�D$P�\$�D$H�$��������ݜ$�   �D$@�\$�D$8�\$�D$0�$���������ݜ$�   �D$p�\$�D$h�\$�D$`�$����������ݜ$�   ݄$�   ���D$8���D$0��݄$�   ������݄$�   �L$@����݄$�   �����L$ �D$����݄$�   �L$(�����D$x���������L$P�D$H����݄$�   �L$X������܌$�   ����ݜ$�   �D$h�����D$`�������D$p�L$@�����������L$ ���L$���D$p�L$(���������D$h�L$P�D$`�L$H���D$p�D$X��������݄$�   �������\$x݄$�   ����݄$�   ������݄$�   �D$@�������������L$ ݄$�   �L$�����L$(�������������L$P݄$�   �D$H���������������������D$x݄$�   ������Az9����������Az\�ٰ����݄$�   �݄$�   �^݄$�   �^^��]� ����������Az#�ٰ�����D$`��D$h�^�D$p�^^��]� �ɰ��^�^^��]� �����V�t$��thH>����A����t��^�3�^���������������̸H>����������̋�P�����������V����_  �N$N��$��^����������̃y ����������̋A��~
�y t���3�������������̋A������������̋A�IPQ��) �����������������̋A(��t�I �L$��� 3�� �����̋A(��t�y t�Q �T$Q��� ��� ������������̋A��t
�L$��� ��� ���������̋D$�QP�A�IRPQ�:) ��� ����VW�|$��F�N�VP�FQRPh =W�-r �N�VQR��( Ph�<W�r �F�N�V��,PQR���| �~ ��<u��<P�FPh�<W��q �F(����uhx<W��q ��_^� �N �Vhp<P�FQ�NRPQ���4y _^� ���������������U������8VW����u �E��th�=P�mq ���e� _^��]ËU��}!�E��tRh�=P�Dq ���<� _^��]Ã�}!�E��tSh�=P�q ���� _^��]ËM;�}"�E��tSQhx=P��p ����� _^��]Å��D$<    ~=3���~!��I �����$���������t%��;�|�D$<�M��;E�D$<�<�|ð_^��]ËE��t���T$<���$VRhH=P�up ���m� _^��]��������U������4SV��V��W'�E��tRh8@P�8p ���0� ��_^[��]� �F��}�M��t�Ph@Q�ϋN;�}(�U��t�PQh�?R��o ����� ��_^[��]� �~ �Bu�V ;Ћ}}��t������PRh�?W�o ���~( u'���j���hx?W�o ���� ��_^[��]� �F��u'���<���hX?W�fo ���^� ��_^[��]� �NWP�FPQ�/ ����u'�������h$?W�)o ���!� ��_^[��]� �V �FWRP��������؋F(�k�������u'�������h ?W��n ����� ��_^[��]� 3�9N��  ��~�����F�V(�L$�E  �F���0'�������������Dz�D$��D$    �F9D$��   �F�������Dz1�������D��   ��������Dz6���������z%���������ʋF ����;ύ�|��������   �������������AzԋE�څ�������������V�ʍʃ��\$�A��$h�>P��m ����� ��_^[��]� �U�څ��������p���Q+ȃ�Qht>R�m ���� ��_^[��]� �E�څ��������7���Qh@>�#����؃~��_�~uY��uT�D$(P���`m  �L$Q����m  �T$R�L$,������t*�E�������h>P�m ���� ��_^[��]� _^�   [��]� ���������̋T$3�9D$��P�D$R�Q(P�A R�QP�A�IRPQ��2 �� ��� ����������j�h�:d�    P��0SUVW�  3�P�D$Dd�    ��\$T3�Uj���gp ��;��e  �FP���j ��;���   �NQ���{j ��;�to�VR���ij ��;�t]�FP���Wj ��;�tKU���Hj ��;�t<U���9j ��;�t-�L$�y# �L$Q�ˉl$P�I� �L$���D$L������# 9nt�N�F;�|��|QP�z" �����tU����i ����t�VRU����i ���F��~�~ t���D$T��D$T    �~( t�D$T��~�n��~9F }3��tLU���}i ����t?��~;3�9~~4��t0�F(��t�N �ύ��3��T$TPR���Vi ��;~��|���ǋL$Dd�    Y_^][��<� �j�h�:d�    PQVW�  3�P�D$d�    ���D$    �|$ ���D$    ������N�V�GP�FWQRP�D$,    �D$    �:* ����u���,����ǋL$d�    Y_^��� �����̃� V��NW3�����  �V;���  9~��  �D$4�D$,��������  �F�D���T$�D���T$��������Dz��������Dz�G��_��^�� � ��������A�T  ����V  �D$4�d$,���D$���D$�������\$����$�\$ �����D$,���D$43Ƀ��D$�D$�D$�D$ ��   �z��F�������F�ȍ�u���������������F�T������F�D��D�u���������������F�T������F�D��D�u���������������F�T������F�D��D�u������������Ń��;��T���;�}-�F�������F�ȍ�u������������Ń��;�|���_�ڸ   ��^�����؃� � ��_^�� � ����_��^�� � ��������������̋A�QP�ARP�O  �������������̋D$�QP�A�IRPQ��  ����� ̋A��|����3�����;S�\$UVW������z��2ۋF�NPQ� �V�N�����i�t	����   �~;���   ����   �~ ��   �~( �   ��u6�~ tu�����un��~%�~��    �\9��������DzP���;V|��D$���   �����$�Ѕ�u+�D$�L$�T$���$QR���U{  ��t_^]�   [� _^]3�[� ������������U����j�h;d�    P��lVW�  3�P�D$xd�    ���Ph�L$4Q��3��ҍL$4��$�   �3�����t`�N�V�D���v�E��������z
�D���\$<��T������Au�D���\$4�E�MPQ���\$�D$\�\$�D$T�$�t�
 �� ���L$4Ǆ$�   �����k �ǋL$xd�    Y_^��]� �����U������4SV��N��W}3�_^[��]� �E ��t� �3��]�E�VP�FS���$PRQ�� �������t��uX�F�E�N�\$8�T$8��D��R���\$�D���$S�;� ����t%�D$8�F�N�U�VWS���$PQR� �����M�E�F �UQ�MR�Ѓ����$Q�N(��R�VP�F���FQ�NRPQ�I �M ��,����t�9_^[��]� ����������V��3�9F~�~|����   �҅�t�   ^Ë�^�#U  ���QSUV��F�N�VWPQR��  �������D$t^�N �~�n(�����׍\� �V���х��l� |8�d$ �F�NUSPQ�q�
 ����t�F ���+�+��y؋D$_^][Y�3�_^][Y������̃�(�D$DP�L$Q�L$4�������������T$���$�D���������  ���D$��������A{~�\$d����A{u�h@�T$l����{�\$l��؍L$,�����$�L$D�����T$�D$l�$������At�������$�������������{!�����T$��������Dz������2���(����������  ��������   �T$d����z��2��0'S�D$`����������uu��������u;�ڍT$0��R�؍L$L������D$���D$�����L$`��������At.��2��������D$x������u*������������������Au�����ذ[��(�����2����݄$�   ��������Au*��������Au�����������������������{�2�������؄�u���u�2�[��(������ذ��(��V3�9qt0�A(��t;�Q �T$�Ѕ�t,�Q�D$�о   �NO  ��^� ���\$����Dz�   �1O  ��^� �����������SV��F(3ۅ�ta�N �L$W�<ȅ�tP�D$� �   �9^~0�@�_�~~�@�_�F��~������R�Gj P�4� ���~ t��N��_���N  ^��[� ����SW���G(3ۅ���   �O �L$V�4ȅ���   9_t[�\$���~0�C�^�~�C�^�G��~������R�Fj P諢 ���O�C��^�ϻ   �"N  _��[� ��L$�Y������D{�q�   �����~E�A���^�~�I�^��؋G��~'������Rj ��V�2� ��^���M  _��[� ��^���M  _��[� ��������������̋A(V3�����   �Q �T$�Ѕ���   9qtX�A��������D{z�A���4D$�����y~�B������X�y~��^�J�X�   � ��^�X�   � ��D$��y��~�B����X�y~���B�X�   ^� �؋�^� ���������VW�|$����|,�F�NPQ�g ��;�}�V�D$�����L  _�^� _2�^� �SV��F�N�VWPQR�Z �N �V���F(P�FQ�NRPQ��
 �� �����QL  ��t��t	_^�   [�_^3�[�����������V���(L  �D$�L$�V(P�F Q�NRPQ�]�
 ����^� ��̋D$�QP�A�IRPQ� ��� ����SV��N$W�|$;��~!�F(��u"��    P�
z�������F(t*�~$_^��[� ��~��    QP�Cz�������F(uىF$_^2�[� ��������������SV��NW�|$;��~G�F��u��    P�y�������~*��    QP��y�������Fu_�F    ^2�[� �~_^��[� ���������������Q�T$2���V���E  �NW�~+�;��3  �~ �)  �~( �  �F��~�~ t	�x�|$��D$����D$    �|$��SU�l$Q�͍�    ��
 ���D$��   �F�E �N�M�V�U�};~ u!�L$����PQ���O����UPR�Ţ ���?3�9~~4�F(��t�L$��V ���3�SPW���F�
 P萢 ����;~|̋|$�F�L$�ȋF�D���\������Au7�v�D���U�E���\$�D���$Q�MRPQW�mP �D$@��$][_^Y� 2�][_^Y� ���̃��Q(��$�$P�A R�QP�A�IRPQ�[ �D$�� ���̃� W��� �|$�M  ��P4UV�ҋo����t$�-  �G ;��"  ���  ;�Su	�^�\$��D$�؋���P���.�������l$ ��   ��F���������������҉D$,�t$$�T$�G(��t�O �͍<��3��L$����|$,�|$�|K�q���T���+��ݍD�����B�� �X(�� ���D �X �B(�X�B �Xu܋l$ �|$�t$$�T$��|�׍�+���������}�T$�D$�|$(�Ã���l$ �t$$�N����\$�؉_ �G   [� ^]��_�� �������̃��|$$ SU�l$4W����t9�|$4 t2��t.��t*��|&�D$$;���������R�L$�v�������D$u	_]3�[���V�t$,���V��u�������D$ u�D$P�v����^_]3�[���Vj U�ݛ �t$ ��3ۃ����L$�\$��   �t$,�D$3Ƀ�|;�V������E��    �@��� �����X��@����X��@����X��@����X�u�;�}�D� ��;����\��|�T$��R�vu���D$$P�lu����^_]�   [��Ët$�L$�\$3�3҃�|o�~��p��;�t�A��l$�\� ���n�;�t�A��l$�\� ��;�t��l$�\� ���n;�t�A�l$�\� ������ ��;�|��l$<�t$�L$;֋|$}��;�t	�у��X���;�|�\$ �L$8�T$4�D$0�t$,SWQ�L$4RPQV�I ������   3���|W�T$,�������+����K�E�<�    ��I �A�� �@؃� ���X��D��@��X��A��@��X��A��@��X�uЋt$,;�}�Ӌ�+ՍD� +�������@��X�u�D$��;D$�D$���������W��s��S��s����^_]3�[����������̃�VW�|$$����}
_2�^��� ;~��  �E  ;~}G�~ ��  3�9N��  �F(��t�V �э��3��V�Ѓ���;N|ۉ~_�^��� �~ S�_u�ߋF ;�}�\$��D$��;�}%�~$ ~�F�N(�ÉF$���PQ�:s�����F(�N���L$�   �������������U�T$�\$$��L$�F(��t�^ �ٍ,��3�~ ��l$ �\$t
�F�D� ���G�;F|�Ã�;F}��N����y��|H�D���T���+\$�����ݍ��B�� �X(�� ���D �X �B(�X�B �Xu܋\$�l$ �T$��|�Ս�+���������}�T$�D$T$$�|$,�����D$�T$�'����\$��]�^ [�~_�^��� ����3��D$����������   �D$�����Aur�����������H'��4��������p@��Az���!����������z�ڍB�������������!������Az������������Au��   ������؋������̋A��~�y t���3��T$R�QR�Q(R�Q R�Q�IRQP�� ��� ������̋A��~�I�@�D���3������������̋D$��|;A�A� �������������V���8A  ��@�@>3�;�t��F�F�F�F�F�F�F �F$�F(��^������Q�D$SUV��W�nUjP蹮
 �~WjP譮
 �NQjP衮
 �^SjP蕮
 �D$H���0��~\�~  ~V�V(��tO�M ��~
�? t���3����3���L$��~*��    �T$�D$WRP�@�
 �N ����;+�D$�<�|܋�FRP�  �NQ��    �D$$RP�
�
 ��_^][Y� ���������������VW���A  �|$��}_2�^� �L$��|��T$;�|�3�9D$�~���N�V�F���Gu��SRQ�F �}
 ��P���R����N �؋F��Q���������u2ۊ�[_^� �SVW���@  �F(3�;�t	9~$t���3ɋF;�t	9~t���3�;ω~�~�~�~�~�~�~ �~$�~(t	Q��n����;�t	S��n����_^[�������̃�W�΋��#@  �G�F�O�ɉN�W�V�G�F�Ft���F � t:�NQR�	 ��P���s����F�NPQ�	 �N��    �GRPQ�A� ���( ��   �V �VR��������F��~�~ t���3��O ����D$�F ;�S�_(�~(u�N�����QSW�� ��[_���U3�9n~5��    ��    �T$�D$�L$QSW诗 |$\$ ����;n|�][_��������VW�|$��;�tW��K  �������_��^� VW�|$W���������>  �~ u+���W`����Dz�Wh����Dz�_p����D{��؋��:����F(�N �VWP�FQ�NRPQ���
 ��_��^� �����j�hH;d�    P��TSUVW�  3�P�D$hd�    �������l$x�D$,P�L$$3�Q�͉|$(�|$4�3U ��;���  �|$ ��  �T$(R�͉|$,�|$(�|$�|$ �|$4�|$8�> ��;�t"�D$$P���> ��;�t�L$Q����= ��9|$}3��;�t�T$R����= ���D$;D$}3��W;�tS�L$0Q���= ��;�t@�T$4R���= ��;�t-�L$8�� �D$8P�͉|$t�r> �L$8���D$p�����^ �L$�T$�D$$Q�L$,RPQ��������u3�;��|$ta�T$R���9= �L$;���}3��Ft�D$�L$PQ� �L$��;�t3��&;�t"Q���n�����;�t�S�D$RP����< ��;��|$t�L$Q����< ���k;�~
9{t���3�;�t���T$R��������9|$~>;�~:;�t:�{ ~.��t0�C(��t�K �ύ��3��L$xPU�}< ��;{��|�3�;�u�������ƋL$hd�    Y_^][��`� �������������U����j�h{;d�    P��(  SVW�  3�P��$8  d�    ��F�N�VjPQR� �����A  �L$,��B �L$|Ǆ$@      ������$�   ������$�   �������$�   �����L$\�����D$,Pj �����������  �V�L$DQ��R����������  �D$D���d$4�T$d�D$T�d$<�T$l�D$\�d$D�T$t�����������������T$|�$� ��������d  ���D$t������A�M  �N��u5���؍L$,Ǆ$@  ������ �   ��$8  d�    Y_^[��]� ��2�ݔ$�   �E��������At�س��;�U�ȿ   ���;�ݜ$�   �����D$\���\$\�D$d���\$d�L$l�\$l�p�����    �D$|PW�������D$|�D$,��ݔ$�   ݄$�   �D$4��ݔ$�   ݄$�   �D$<��ݔ$�   ���d$Dݔ$�   ���d$Lݔ$�   ���d$Tݔ$�   ����������������������������������������u<���������L$d���L$\��݄$�   �L$l���T$t��A������A��  ���7�����L$\�������L$d�����L$l�����T$t��A��������  �Ʉ������D$,�����L$D��ݔ$�   ���L$4���L$L��ݔ$�   ���L$<���L$T��ݔ$�   t6�܍�$�   Q�؍�$�   ��R��j ��j��
 �����/  �D$t���^�D$|������݄$�   ����������A��   ݄$�   ��������������������   ݄$�   ��������������A��   ݄$�   ������z!������z��������Au�����ݔ$�   ������Az#��������Az�؋V����;�������'������؃���$�   �$P�L$8��? � �\$|�L$|�@Qݜ$�   ��$�   �@ݜ$�   �����]����Az������������������������؍L$,Ǆ$@  ����� 3���$8  d�    Y_^[��]� ���U����j�h�;d�    P��(  SVW�  3�P��$8  d�    ��   9~u*�E�E���$P�s  ��$8  d�    Y_^[��]� 3ۍL$t�\$@�Y�����$�   �M�����Rh��$t  P����S�ȉ�$D  ������ SS��$�   Q��$�   R�����$�J  �����$t  ��$@  � �E����   �����$�҅���   �}��tn��$t  P����I  P�L$xQ��$�  ��  �E���$W��$�  Ǆ$L     ��@ ��u����$��$�  W��@ ��$�  ��$@  � �D$@   �  �~�  ��$�   �1� ��$�   ��$@  �.�����$�   �"����L$\�����L$D�����$�   �\$,�T$|�D$t��$�   �L$x�\$l��$�   �T$d�T$L��$�   �D$\�\$p�D$D�\$X�^�T$T�Ù��?|$h�|$P�������L$`�L$H}�   ���D$(   �S  �L$(��$�   PQ���s����T$(�:;É�$�   �D$(�  �L$(��$�   PQ���E����T$tR��$�   P��$�   �,���P�L$xQ��$|  R��$�   ����P��$�  P�������������D$,��������   ��$�   �\$,��$�   ��$�   �L$\��$�   �T$`��$�   �D$d��$�   �L$h��$�   �T$l��$�   �D$p��$�   �L$D��$�   �T$H��$�   �D$L��$�   �L$P�T$T�D$X��؋D$(�;F�D$(�������$�   �^;ÉD$(������L$DQ�T$`R�D$|P��$   �ً ����  ��$$  Q��$�   �-�������$  �$R��$�   �������L$<�$�����L$,�[������8  �D$4������4��������u-�������T$,����Az���\$,�T$4�@�0'�\$,�T$4�0�D$,��������Az!����������Az����0'�T$4���\$,��$  ��$  ��$  ��$�   ��$  ��$�   ��$$  ��$�   ��$  ��$�   ��$0  ��$�   ��$(  ��$�   ��$   ��$�   ��$�   ��$4  ��$�   ��$�   ��$,  P��$�   ����$�   �$��$D  ��$�  Q��$�   �*����D$<��P��$x  R��$�   P����$�  �$Q����������%����D$4���$  �H��$  �P��$  �H��$  �P��$�   Q��$   �@����$�  �$R��$0  蛷���D$<��P��$�  P��$�   Q����$   �$R�p��������ƶ�����$$  �P��$(  �H��$,  �P��$0  �H��$4  �P��$8  �E����   ����$�   �$Q���҅��D$@t�}��t�    ��$�   󥍌$�   Ǆ$@  ������� �D$@��$8  d�    Y_^[��]� �������������̃�SV�ً�PWj �ҍL$�������3���t:U�l$,;s}/�D$PV��������L$Q��軆 ���\$0����Au3�����u�]��_^[��� ����������D$4����A������z�������A������z?��������Au�������0'�(���������%�$��������u	������At�������A�L$�T$ ��@�\$8���5���\$H��&�\$@݄$�   �\$8�\$0��L$|�P��$�   �H��$�   �P��$�   �H�L$\�P�T$`�ĉ�L$d�P�T$h�H�L$l�P�T$p�H�P������X�����������L$�T$ ��@�\$8���5���\$H��&�\$@݄$�   �\$8���\$0��L$|�P��$�   �H��$�   �P��$�   �H�L$\�P�T$`�ĉ�L$d�P�T$h�H�L$l�P�T$p�H�P������X�����Ã� VW���P3�W�҅���   �D$,P�L$Q���VA  ����������   �F��~
9~t���3��V�N(jR�V Q�NR�VQRP�h ����T$9~t$�F(��t�N���ȃ��T$�L$4�$�x�����؍T$,Rj ������9~t�D$���$j ���>������-  _�   ^�� � ��_^�� � �� SV���Pj 2��҅���   �D$,P�L$Q����@  ���.�������   �F��~�~ t���3��V�N(jR�V Q�NR�VQRP� ����T$�~ t.�F(��t�N�؃��N N�ȃ��T$�L$4�$英����؋F�T$,R��P��������~ t�N�D$�����$Q���F������,  �^��[�� � ^��[�� � �������U����j�h<d�    P��   SVW�  3�P��$�   d�    ��F�N�VPQR��
 �؃�����  ��Pj ���҅���  �L$d�b9 ��P0j��Ǆ$�       �ҋF��~�~ t���3��N�V(jQ�N R�VQ�NRQP�< ����u.�L$dǄ$�   ������: 2���$�   d�    Y_^[��]� ��Bx���ЋN�����_��Q�Ή|$T�$����V���׃��V R������S�L$h�9 ��D$`P�B|���ЋF3�;�~9^t���D$X��\$X3ɋǺ   �������3��������P�U@�����D$\;�Ƅ$�   th�h��W�XjS�8详 �N�\$T�^����;�Ƅ$�    �D$\    ��   �T$T���T$L9|$\��   �F�D��������A��   �V�F�L$LR�VP���R�>�
 3�9~~3�F(��t��+N�T�V ���3��L$LPjW����ܧ
 ��;~|͋F�D��|$L���\$��+N���$�T��G�R�W�P�D$pQRP��0 ��$�   ��$���|$L�|$P�N����;��/����V���׃�3�9|$P�V��   �L$`�D$T�L$X�D$\3�9^~n�L$\S��
 �N�V(����˅҉D$LtB��|>;N}9�F ���N�ɍ�~�~ t���3ɋD$L���QPR�� �����b)  ��;^|��L$X�V��3���~ �V��^����Ѓ��ӋV��;�|��D$\����;|$P�L$X�F����N��3���~'�L$`�V���^���T$PЃ��ӋV��;�|݋D$T��t�H��x�h�QjP�� W�,?�����L$d�Ǆ$�   �����7 �} �,  3�9~�!  �L$l��
 �V�F�N�T$l�V �D$p�F(�L$tW�L$pǄ$�      �T$|��$�   蚥
 ��$����D{F��P0j���ҋF;Fu������P�L$p�i�
 �F���$����P���$W��$�   �w�
 �F(;�t�N+N�N �ȉT$|��|$|�F��P�L$p��
 ��$����D{7��B0j����W�L$p���
 ��N���$��Q���$W��$�   ��
 �L$l�|$|Ǆ$�   ������
 �Ë�$�   d�    Y_^[��]� ���j�h8<d�    P��(SUVW�  3�P�D$<d�    �����   �ҋ��Ph�L$,Q�Ήl$��3ۍL$,�\$D�Z������L$,u�D$D������� �  S����� j�\$ �L$0�	���� �L$,�\$$�D$D������� �|$T���R  ;��J  �D$�D$L�������  �D$$�������  ��������Dz2;�����uS�������"  ����  h�Bh�Bh�  ��  ������Dz/;�uj���d�����  ����  h8Bh�Bh�  �  ����%  ��~����   ���҉D$T��\$T�D$L�F�N�VSS���$PQR��
 �؋F��F ��P�Ή\$ ��������j  ���z����P��� ������Q  �V�F(�L$Q�N R�VP�FQRP�Ή\$0�����D$dPW���$�3 ��(��~F�|$T ��   ����   ���Ѕ���   �N�V�FQRP���
 ������   �~3�+�����   ��l$�E�9D$��}#S�������F(��tT��|P;~}K�N �ύ��!W�������F(��t1��|-;^}(�V �ӍЋ��S������PUR�} �����$  ����;\$|���Fj��������9�������h B��h�Bh�  �h�Ah�Bh~  hx@�
� ��2��L$<d�    Y_^][��4� ���������������U����j�hh<d�    P��hSVW�  3�P�D$xd�    ��]���8������?  �F��~�~ t���D$��D$    ��~�Ph�L$4Q�Ή|$$��P��Ǆ$�       �Z����L$4��Ǆ$�   ������ ���c  ���e#  �E�@�N�V�T$$j j����$QRW�3�
 �D$@�N�\$H�؍;�D�����\$�D���L$<�$��������t �F�D$,Sj����$P�FPW���
 ���؋F(��t�N �ˍ��3��D$$�V���\$����V �$j�QP�D$8RWP�T! ��(��u3h�Bh�Bhl
  hx@�d� ��3��L$xd�    Y_^[��]� �;PW�F��
 �N������;�|�D$$�V�N����;�}��؋U��F�N�T$$j j���$PQW��
 �D$@�N�\$H�؍;�D�����\$�D���L$<�$��������t �D$,�F�VSj���$PRW���
 ���؋F(��t�N �ˍ��3��D$$�V���\$����V �$jQP�D$8RWP�4  ��(��u3h�Bh�Bh�
  hx@�D� ��3��L$xd�    Y_^[��]� �N��+�;��D$��   �F ��������+�3Ƀ�|8��V(���ʋV(�D����\��V(�D���\���V(�D���\���W�;�|�;�}��    �N(�������;�|�F�L$ PQ�}�
 ��+���3҃���|7�X��~�σ��׋~�D���;��\��~�D���\���~�D���\��|�;�}�<�    �V�ʃ��:��;�|�T$�|$ �V3����x�D$$�N����;�~��؋F��~�~ t���3��V�N(jR�V Q�NR�VQRP�c�
 �����	   �   �L$xd�    Y_^[��]� ���������������U����j�h�<d�    P��hSVW�  3�P�D$xd�    �����   �҅�t2��L$xd�    Y_^[��]� �3�9F�������B4�Ћ�RhǉD$�D$$P���D$ ��j ��Ǆ$�       荛���]j �ˋ�菛����D$����{�D$ �L$$Ǆ$�   �����(� �|$ ��   �F��~�~ t���3��N�V(j Q�N R�VQ�NRQP�-�
 �V�~(��j �ˉT$�����F�N �T$���\$���$jP�D$4WQRP�A �F�����(3���~��j ���ך���N���F�����;�|��D$��Rh�D$4P����j��Ǆ$�      荚��j�ˋ�蒚����D$����At�D$ �L$4Ǆ$�   �����+� �|$ ��   �F��~�~ t���3��N�V(jQ�N R�VQ�NRQP�0�
 �F�~+��D$<�F(����t�V �׍ЉD$��D$    j��������N�D$���\$����N �$j�R�T$8P�D$8QRP� �N�VQR� �
 ���F������0;�|j��襙���N���V����;�}��D$��|$ t���-  �D$�L$xd�    Y_^[��]� ����j�h�<d�    P�� SUVW�  3�P�D$4d�    ���D$L����D$(    thH>��������T  �L$P�	��thH>��������8  ��Bj ���Ѕ���  �O�W�D���D$D��������A��  �G�\��������  �L$L�1�T$P������u/j,�{0�����D$,���t$<t��������l$<���3��l$<���;���  ��u+j,�@0�����D$,���D$<   t	�������3��l$<�؋���  ����  �D$D�G�O�Wj j���$PQR��
 �D$`�O�\$H��G��D�����\$�l$,�D���L$<�$�.����D$<����tH�G�O�T������A��   �W�T��������   �GUj���$QRP�8�
 �D$H����D$���S  �W�G��+�;��A  ���ʺ���Oͅ�D$�L$��   �W�A��D$,����D$(����D��  3�;O|y�D$(�D$ ;T$,��  �D$ � ������DzT�l$ ����;O}׋W�؉L$�B�L$L�؃9 u��t��Bj���ЋL$P�9 u��t��Bj����3��  �L$�W�؋G+�;ȉT$ �2  ;��*  ;�t�G�F�G�F�G�N�L$�F�N ;�t�G�C�O�K�G�L$�C�S�K �V(;W(tY�D$�D$P������3�9l$~@�l$$��D$���PU���͹���N(L$(PQ�?r �D$ ���D$0����;l$|ŋV;Wt3�D$�OPQ�?�
 ����U�������G�N��    RPQ��q ���S(;W(u�|$ ~|�l$ ���D$P���h���3�;�D$$~_�D$(�G(��t!�L$�T$$��W ����L$�W������3��l$���UP�C(D$0P��m �D$0l$4����;D$ �D$$|��K;Ou�|$ ~:�T$ �GRP�r�
 ����U���E����W�D$��    Q�SQR�m ��;�u�D$ �L$�C�K ;�u�T$�D$�V�F �F�N(+F��t�V �Ѝ��3��D$D�V���\$�����$j�P�D$,Q�OPQP�� �F�VPR�h����
 ��0;�})���    �F�D$D��N�VQR����
 ��;�|ߋF��~�~ t���3��N�V(jQ�N R�VQ�NRQP��
 �D$`�S�\$��C(�O�\$��jRP�D$0PQP�5 �S��(3���x�D$D�K���S����;�~��؋C��~�{ t���3��K�S(jQ�K R�SQ�KRQP��
 �D$h���8 u�0�D$P�8 u��D$(   �>�T$L�: u��t��Pj���ҋD$P�8 ��������������Bj����3���؋D$(�L$4d�    Y_^][��,� ����V�t$W���   �~����D$��t�P���   ���Ѕ�u_^� ��_^� ���������j�h=d�    PQVW�  3�P�D$d�    j,�*�������t$3�;��|$tG���<  ��@�@>;�t��~�~�~�~�~�~�~ �~$�~(�ƋL$d�    Y_^���3��L$d�    Y_^�����������j�h;=d�    PQSVW�  3�P�D$d�    ��j,��)�������t$3�;��|$t5���  ��@�@>;�t��~�~�~�~�~�~�~ �~$�~(�3�;��D$����t;�tS���Q"  �������ƋL$d�    Y_^[��������VW�|$��t@hH>���:�����t0�t$��t(hH>���"�����t;�tW����!  ������_�^�_2�^��j�hh=d�    PQVW�  3�P�D$d�    ��t$�  3���@�@>;ȉD$t��|$ ;��F�F�F�F�F�F�F �F$�F(tW���o!  ���8����ƋL$d�    Y_^��� ��j�h�=d�    PQV�  3�P�D$d�    ��t$�#  3���@�@>;ȉD$t��L$$�T$ �F�F�F�F�F�F�F �F$�F(�D$(P�D$ QRP�������ƋL$d�    Y^��� j�h�=d�    PQV�  3�P�D$d�    ��t$��@�D$    ��������D$�����  �L$d�    Y^��������U����j�h >d�    P��XSVW�  3�P�D$hd�    ��V�L$<�H����D$T�L$L�T$HPQR�D$|    ���
 �L$T���D$XPQ�|$8��
 �L$\�D8��+����F�D$`3҃�3����N�T$~{��T$�L$T��t�����R�\$0�T$LQPR�h�
 �؃���|:�C�D$ ��|%�N�VQR�7�
 ��;�}�F�D$,�����o  ���l$ u͋L$�D$L�;ȉL$|��N$�V(���Q3�SR�f �~��;�~9^t���|$��\$���D$$3Ʌ��\$�L$ �  �D$$��I �L$ �\$�F�؋D$T�T$,�ȋD$`3�;ǉT$(t�T$X�эЉD$��|$�F(;�t	�N �ˍ<ȋ���   ���ЋN�V�D�P�FQRP�S�
 �N�V ��+��Ӄ�;ٍ<�}6�D$(�L$�T$XWP�D$ Q�L$TRPQ�L$D���W����V ����;^�<�|ʋT$�F�NR�VRPQ���
 �L$d�T$\�D$,�D$0P�D$\QRP��
 �� �l$$�D$ �����|$�\$`�V(3����\$�T$(�D$|T�K+ڍB�W����\$,����    �\$�\$,�A�� �X؃� ���D��X��A��X��A��X�u܋T$(�\$�D$;�}��+�+L$��������X�u�D$`3�;�t�L$L����L$X�ȉT$��\$�V(;ӋFt����F ���3҃��T$$|H�t$�L$�B+�W���������    �A�� �X؃� ���D��X��A��X��A��X�u܋T$$;�} �L$+ʍ�+���$    ������X�u��D$8�@�L$8�D$p   �  �D$`3�;�t9t$\u3��|$T;�t9t$Pu3�;Ɖt$@�t$D�t$H�t$L�t$P�t$T�t$X�t$\�t$`t	P��=����;�t	W��=�����L$8�D$p�����x  �   �L$hd�    Y_^[��]�VW�|$����|�F���;�|u_�^� j�9�����u_2�^� ����   SU���ҋ+��F�D$�Bx�΋��ЋN�VQR���m�
 ��������W���8�����t?+|$��+����~ W������t&3���~��I ��������t��;�|�][_�^� ][_2�^� ������������U����j�h(>d�    P��`SVW�  3�P�D$pd�    ��~ �}�D$ u6;�tW�
  ���������Pj ���҅����L$pd�    Y_^[��]� � t�~ u�]�������  ����   ���ҋ؋���   ����;�~����   ����P���s������b  ��P4���ҋ؋�P4����;�~��P4�����P�Ct���Є��/  �~ t
� ��  ����   ���Ћ�؋��   ����;���  �O�W�Gj QRP���
 ������  ��B4���Ћ�؋B4����;���  ��Bj ���Ѕ��Z  ��Bj ���Ѕ��G  ����   ���Ћ�؋��   ����;��%  �~ ��� ��:��  ��P4���ҋ؋�P4����;���  j���������8  j ���x����\$$�^�C�P���f�����~ �\$,t���D$$��������D{���\$,����؋O��N Q���,����F�O�V�QR��
 ��P�������F�P�R���1����\$$�G��P�������l$$R���\$8迫���΋��f����O�L$$�ωD$脫���ΉD$ �y����W��;T$ }3����D$�I R���ȫ���D$4�D$�N�����;T$ �D$|ڸ   9D$$�D$��   �D$�V ���P�D$ P�ύ��*���PS�c ���D$8����������D{^�T$3Ƀ�|?��������C��    �@��� �����X����H��X��@����X��@����X�u؋T$;�}�˃�;����\��|��D$�؃F��;D$$�D$�O�����L$pd�    Y_^[��]� �D$�L$pd�    Y_^[��]� W�L$D�|�������   ���D$x    ��P�L$D������u(�L$@�D$x�����i���2��L$pd�    Y_^[��]� ��B4����P�L$D������t��~ t�L$@�|�����t�j �L$D������t��~ ���|$L ��:�u��D$P��|�x��3�����   ����;��h�����P4�|$H����;��L$@t$�D$x���������2��L$pd�    Y_^[��]� j �b������ ����D$@P��������L$@���D$x�����{����ËL$pd�    Y_^[��]� ����V��F�V;�u?�@��Ɂ�   v��|�]UU ;�}�������   ��;�}P���k���N3��I�N�щ�A�A�A�A�A�N�F�I���N��^��V��������D$t	V�������^� ��U����j�hn>d�    P���   SVW�  3�P��$�   d�    �����   �҅���  ��Ph�L$\Q�����E���T$\�L$d�$Ǆ$      諄������������At	������z+�v ��������Au��$���L$d�$�0����\$T������D$T���L$d�$�S������D$T�   S���L$h�$�8������  ��$�   �D����L$l��$   �4����D$T����   ��$�   �D$P�L$l�L$L�D$LP�L$TQ�����$Ƅ$  �ҋ���t,��$�   P�L$p������L$l;�t��R���  �D$l������L$l��$   �7�����$�   Ƅ$    �#�����t#��L$\�����E�Cl�����ɋ��\$�$�ЍL$\Ǆ$   ������ �ǋ�$�   d�    Y_^[��]� �������������U����j�h�>d�    P���   SVW�  3�P��$�   d�    ��]3�;؉D$,t9C|�C�};�t9G|�G�P�B�Ѕ���  �F��u|�ۋF�D$,t09C}P����h��3�9~~��������PW���P�����;~|�}����  �F9G}P����i��3�9~��  ���N���MR�������;~|��b  �\  �N���P  ���G  �^�~+؃��L$<�|$8�\$l�m �L$|Ǆ$       蹈����$�   譈���D$TPj ��蟷��3ɅۉL$0��  ��F�D���\������A��  �^�D�������D�+  �Ë����D:��\������D�  �D$T�T$X�D$<�D$\�D$D�D$d�T$@�T$`�D$L�D$TP�L��T$L�T$lQ�ΉT$X�����   ���;߉|$4�@  ��$    �D$0�T$|�RQ���ܶ����T$t�\$tR��$�   P�L$D�  ���}  �N���L$p�D$p�L$<�D$t���D$4�������p&����A�  ����$�   �$R�� � ݔ$�   �@ݔ$�   �@ݔ$�   �D$|�����������������P+����;������������A��  ݄$�   ������������������������������  ݄$�   ����������������������������A��  �F����;��|$4������D$,�|$8�\$l�L$0����;ˉL$0�|$8� ����|$, ��   �}�D$,��u	9}��   �L$|Qj ���b�����t�T$,R����m��������Pj ���A����}��t�D$,P�������N�V�D��P��������~�D$0    �F�D���\������Au4�M��t�c����N�T$0P�D
�P���ߴ���M��t�V�D��P�����D$0����;ÉD$0|��L$<Ǆ$   �����E� �]����   ���Ѕ���   �|$,��   ����   �C��~g�K�d��Ǆ$   ������� 3���$�   d�    Y_^[��]� �������؍L$<Ǆ$   ������� 3���$�   d�    Y_^[��]� 3Ʌ�~�@�C�D���3����Q�P�Q�P�Q�P�Q�P�I�H�D$,��$�   d�    Y_^[��]� �����������V�t$��th8?���K�����t��^�3�^���������������̸8?�����������V���h1
 ��C��^��������������̋D$VP���c1
 ��C��^� ���������C�1
 ���������������������j�h�>d�    P��V�  3�P�D$d�    ��@h�T$R3��ЍL$�t$ ��}����t+�t$(��t�L$茑����t$,��t�L$������   �L$�D$ �����1� �ƋL$d�    Y^��� �����������̋�P0j���������j�h�>d�    PSVW�  3�P�D$d�    ��L$ �D$    �}����t7�>j�L$$��{��j �L$$����{������\$��� �Gl�$�Ѕ�t��2ۍL$ �D$�����|� �ËL$d�    Y_^[��� �����V�t$��~��P4��;�u	�   ^� 3�^� �������������SV���PxW3��ҋ�����   ��   P�K-����؋B|��S���Ћ���tc�L$�D$j Q���$S�WRj��
 ����|=;�9�L$��t��L$ ��t)�D����\$���$趌��S� -����_��^[� 3�S�-����_��^[� _^��[� ����������j�h(?d�    P��V�  3�P�D$d�    ��@h�T$R3��ЍL$�t$ �{����tBj�L$�Rz��j �L$���Ez���D$(�L$4�T$0QR���\$��\$� �$���
 �� ���L$�D$ ������� �ƋL$d�    Y^��� �����j�h[?d�    P��   SVW�  3�P��$�   d�    ��L$� ݄$�   ���$�   ���   ���$�L$QR��Ǆ$�       �Ѕ��Ä�t+��$�   ��t ݄$�   �    �t$ݐ�   ��ݘ�   �L$Ǆ$�   �����p �Ë�$�   d�    Y_^[�Ĥ   � ���U����j�h�?d�    P���   SUVW�  3�P��$�   d�    ����P42ۈ\$K�ҋ�����  ��Ph�L$TQ���҃�Ǆ$       ~����P�*�����D$L�
�L$d�L$L�����j jPV��j ���,��$�L$p�l� �T$l�x���D$d���   �����$�҅��!  ���j j�UVj ���L$p�$�D$l�Sx���T$d���   �����$�Ѕ���   �L$LUQj V虣
 ������   ��pDj j SVj ���L$p�$�T$l��w���D$d���   �����$�҅���   ��hDj j �D$X��PVj ���L$p�$�w���T$d���   �����$�Ѕ�tP�L$LSQj V��
 ����u;�<�WUj V��
 ����u'SUj V�ޢ
 ����uWUj V�͢
 ����u�D$K��~�D$L��t	P�n)�����L$TǄ$   ������� �D$K��$�   d�    Y_^][��]��Ë�$�   d�    Y_^][��]��3�� ����������́�   SUV���P4W�҃���$  ����U �U�]�0��P4����=�   �|$���P4�������P�w(��������$$  ��$   ��S4PQW����݄$   P���   j �����$�Ћ�؋B4���Ѓ�~*���B4�] �G���]�G�]��=�   ~	W�G(����_^]��[��   � �����2�� �����������U������4  ��P4SVW�L$<����]��S����@�S�E��P�X�|$@�����P�'�������E�E�L$<����   P�EPWVj���$�҃���M����D$<�~1���G�[�D��Y~��@�G�[�D��Y~W�o'���D$@��_^[��]� ���������������U������4  ��P4SVW�L$<����]��S����@�S�E��P�P�E��P�X�|$@��v���P�&�������E �E�L$<����   P�EPWVj���$����U�D$<�����������8�8�E�~9���G�[�D��Z�A�X~!��@�G�[�D��Z�A�X~	W�t&�����D$<_^[��]� ����U����j�h�?d�    P���   SVW�  3�P��$�   d�    ���G��|3��.�u���u@�O�w+�yFh�Dh�Dh�  h�D�4g ��2���$�   d�    Y_^[��]� ��|ƋO�G+�;���W�2�W�D���\������Ath�Dh�Dh�  렋���D��������Dz��G�ʍ0�F�D���\������Dz��L$|�Iz���L$d�@z���L$4���
 �O�T$4R�\1�V��Ǆ$      ��������  �D$LPS���������L$4uǄ$   ������ ������
 �]�����Q  ���;��T$$�\$,��   �L$|QV��豨�����L$4t��T$$R��$�   P���
 ���  �D$$�T$,����A��   �xD��������   ����$�   �$Q�L$@���
 ��T$d�H�L$h�P�T$l�H�L$p�P�T$t�@�L$dQ��$�   Rj j��$�   �p�
 ����u2�D$$����$�   �$P�L$@�^�
 P��$�   �q����]����AzU�D$$��;��\$,�����}��t�   �t$4�L$4Ǆ$   �����>� ���$�   d�    Y_^[��]� �؍L$4Ǆ$   ������ �������������2�� �����������j�h�?d�    PSVW�  3�P�D$d�    �ً|$ ����u+j,�������D$ ���|$t	���T����3��D$�������L$,�D$$����   Q���$V���҅�u*��u��t��Pj����3��L$d�    Y_^[��� �ƋL$d�    Y_^[��� ����̋D$�D$�3�� �VW�|$��;~t_S3�;�~>9~~�~�N��PWQ����;ÉFt4�N;�~��+�R�SQ�:H ��[�~_^� �F;�t�SP�B�Љ^�^�^[_^� ��������������̋Q��t�A��~��Pj R��G ���̋A��    ��   v��|�  ;�}���Ã��   ����������������V����C��#
 �D$t	V�E	������^� ������������VW�|$��;�t��P0j��W���#
 _��^� ������������U����j�h@d�    P��h  SVW�  3�P��$x  d�    ��}$���D$@ t�    �E�]����D��  �E2ۃ�����\$B�\$A�\$C��  �$��N����\$B�
�D$C�D$A��Ph�L$DQ����j�L$HǄ$�      �[n��� �]����Auj�L$H�Dn��� �]����Azj�0j �L$H�)n��� �]����z'j �L$H�n��� �]����uj �L$H��m��� �]j�L$H��m��� �]����Auj�L$H��m��� �]����A{6j �L$H�m��� �]������  j �L$H�m��� �]������  ����   ���҅��U  ��u
8\$A�b  �L$l�t����$�   �t����$�   �t����$�   �st����$  �gt����$�   �[t��j �L$H� m��� j j��$  Q��$  R�L$|Q�����$���������  j�L$H��l��� j j���$�   R��$�   Q��$�   R�����$��������  �ۋD$l�L$p�T$t��$�   �D$x��$�   �L$|��$�   ��$�   ��$�   ��$�   ��$�   ��   ��$�   �y����4����$�   �$P��$�   Q��$  �au������{����u��t�   �E�U��D$@��  �|$B ��  ��$�   �Cy����4����$�   �$P��$�   Q��$$  ��t�����{������  ��t�   �E�U��D$@�  �|$A ��  ��$�   �r����$,  �r����$�   �r���L$T�r����$�   P��$�   Q��$  R��$  P�ӆ
 �L$dQ��$@  R��$�   P��$�   Q豆
 �� ��$,  R��$�   �jt���E(��������Au����t�   �E�E��D$@��   �|$C ��   �E0�L$T�T$X��(�\$ �ă��\$0���$�   �P��$�   �H��$�   �P��$�   �H��$�   �P��$�   �ĉ��$�   �P��$�   �H��$�   �P��$�   �H�P�ٽ����@��u4��t�   �E�E��D$@���t�    �E�M��D$@��؍L$DǄ$�  �����ʸ �D$@��$x  d�    Y_^[��]�0 ���I�I�I�I�I����������V�t$W���T$���T$���$�q���D$j j V�����$�������u3��������N����V����F����N����V_��^� �������������j�hH@d�    P��VW�  3�P�D$d�    ���Ph�L$Q���ҋ��D$$    ��}���|$,���$W���*����L$�D$$����詷 �ǋL$d�    Y_^��� ���j�hx@d�    P��VW�  3�P�D$d�    ���Ph�L$Q���ҋ��D$$    ��}���|$,���$W�������L$�D$$�����)� �ǋL$d�    Y_^��� ���U����j�h�@d�    P���   SVW�  3�P��$�   d�    ��$�   �0o���L$L�'o���}���q���E�]�E�MSPWQ�����$� ������D$��  ���Mv������  �M�ES�]S�T$TR��$�   PQ�����$��������  �T$L�D$P�L$T��T$X�G�D$\�O�L$`�W�G�O����u�������D$�U  ��Rh�D$,P�������T$<�L$,�\$DǄ$       �<h�����  ��E���   �L$DQ�T$@R�����$�Ѕ���  ��$�   �n���L$|�n���L$d��m����j�\$(�L$0�f��� �E��������z��}��j �L$0�f��� �E��������DzM�D$D���T$$��������t/�����L$4�\$��'�$�}f���\$������   �B  �����9  ��j �L$0�3f��� �E��������Au��|��j�L$0�f��� �E��������DzB�D$<���T$$��������A{������L$4�\$��D�$��e���\$����A��   �E�D$$3ۉ\$ �\$��E������������D{{�Mj Q�T$lR��$�   P��$�   Q�����$�v�����tQ�T$dR��$�   ��n����������{1������Au�D$ ��D$�D$$������$�T$$�w�������؋D$ ��~�L$ȃ�u���ws���L$,Ǆ$   �����ó �D$��$�   d�    Y_^[��]� ������̃�0V��L$��k���L$��k���D$8�D$P�L$LPQ�L$H�T$R�D$(PQ�����$������^t�T$D�D$@RP�L$Q�T$$R� �
 ����0� �������U������4SVW��W�<�������t&�M�EQ���\$���E�$j ����_^[��]� W��
 ������t{���Y	 �������C  �U���8  �N�9�:�y�z�y�z�y�z�y�z�I�J�N�q���r�q���r�q�r�q�r�q�r�I�J_^[��]� W�ߑ	 ����t�}��t
�p�   �_^[��]� W�� ����t5j ���F- ����   �U�ER���\$���E�$�����_^[��]� W�$�	 ������ta���� ����tT���w�	 �E�uV�����\$�E�D$S�$��t������=   �؄�t�|$? t��t�����
 ��_^[��]� 2�_^[��]� ���������������U������4SVW��W�|�������t+�M�E�P+PQ���\$���E�$R�S���_^[��]� W�4	 ��������   ��� ��|b�M��t[�~�T@��׋:�9�z�y�z�y�z�y�z�y�R�Q�v���@�T��2�1�r�q�r�q�r�q�r�q�R�Q3Ƀ�����_^[��]� W��	 ����t�}��t
�p�   �_^[��]� W�� ������t>��������P���l+ ����   �U�ER���\$���E�$����_^[��]� W�J�	 ������ta���:� ����tT��蝫	 �E�uV�����\$�E�D$S�$��t�j���������؄�t�|$? t��t����
 ��_^[��]� _^2�[��]� ������D$�D$j ���\$�D$�$P����� ���������������V��~ ��Dt%�F��tj P��D�F    �F    �F    ^�����������VW���w��~3��I �G���<� ��t� ��t��ȋBj�ЋO��    ��ҋG��t�W��Rj P�;8 ���G    _^���������������UV�t$j ��h � @���ڕ ��tyj j���k� ��tj�ESWP���� ��3���t?��;}}8�E�<� ��tj�y� �؄�t�M��R���� �j �\� �؃���uË��< ��u_[^]� _��[^]� �������̃�UV3�W���t$�t$�t$�t$ �t$$������l$,�D$ P�L$Q���8+ ���  �|$ � @S������   �T$ R�D$P���� ����   �|$��   �L$0Q���� �؄���   �T$0R����  �D$0;�|;G�G�������;t$0}v��tr�D$P���D$     �a� �؄�tM�|$uF�L$Q���D$    �`� �T$��R��������O���W���<� u�L$��t	��Pj�҃���u��2ۋ��|  ��u
[_^]��� ��[_^]��� ��V��~ ��$t%�F��tj P��$�F    �F    �F    ^�����������U����j�h�@d�    P��hSVW�  3�P�D$xd�    �E�p��Rh�D$4P2��҃��}Ǆ$�       ������`  �E���$�]�������G  �]�{ ~�C�3��E���$VP�*z
 �����|�N�;��S���]����Dz��2ۀ} ��   ����   j�L$8��\��j �L$8�D$4��\���L$0������\$� ���$��
 ��M����|e�V�;�}^�U�B�D���� ��$�E������z�B���$�������Az�س���k��������Au^�R�l�������AzR�����I;�u�E�E�H�d��������Az/�����7�&��} �U�B� �e������Az��    ����؍L$4Ǆ$�   ����迪 �ËL$xd�    Y_^[��]� �������̋D$V��3�;���D�N�N�N~P����  ��^� �����̋D$V��3�;��%�N�N�N~P���\C����^� ������V��~ ��Dt%�F��tj P��D�F    �F    �F    �D$t	V��������^� ������U����j�h!Ad�    P��(  SVW�  3�P��$8  d�    ��]��t�M�mn����u
3ۋM诩 �D$DP�������}��t=�L$DQ��$�   R��������L$D�P�T$H�H�L$L�P�T$P�H�L$T�P�T$XS�]�D$HP���� ��$�   Q����������T$D�H�L$H�P�T$L�H�L$P�P�T$T�@�D$Xt=�L$DQ��$�   R���������L$D�P�T$H�H�L$L�P�T$P�H�L$T�P�T$Xj�D$HP��蘯 ��$�   Q����
 W��$�   RSǄ$L      ��S
 ������   �L$`�+��������   j ���L$l�$Q��Ƅ$P  �҅���   �D$p����   9D$t��   ��$�   �R
 �L$t�D$p3�+�Ƅ$@  xS��$    �L$|��D���\������Au&��$�   RV�L$h�ّ����tWjS��$�   �%R
 �L$t�D$p��+�;�~���$�   Ƅ$@  �P`
 �L$`Ƅ$@   �������$�   Ǆ$@  ����舧 ���$8  d�    Y_^[��]� �L$`Ƅ$@   ������$�   Ǆ$@  �����F� 2���$8  d�    Y_^[��]� ������������U����j�hqAd�    P��(  SVW�  3�P��$8  d�    ���|$H��P43��҃�t��P4���҃���  ��Px���ҋ�����   �ωt$D�҅��D$,��  3���;��D$4%�D$8�D$<�D$@~V�L$8�?��3�;���$@  |
;t$@�t$<�L$8��P|Q���҅���  ���]����Dz	��;�]��$�   P������P��$�   Q���	���P��$�   謥 ��$�   Ƅ$@  �x�
 �]����A��  �L$|�W����L$L�\$dƄ$@  �   �%^��3�9|$D�E  �T$,�D�D$0�D$0�����\$t�D$8�D����\$��$�   ���$�h��3Ʌ�����;t$0�L$,��   ���$    �D$,����$�   �L$|�$�V���L$H����$�   �$R������L$L�P�T$P�H�L$T�P�T$X�H�L$\�P�D$lP�L$PQ��$�   �T$h��
 �D$l��t�D$d������At�xD������z3ۃ���$�   �$R��$�   ��
 P�L$P�t���]����Au3��D$l��;t$0�\$d�t$,�!�����;|$D������L$|Ƅ$@  �c� ��$�   Ƅ$@   �O� �|$@ Ǆ$@  �����D$4%t�D$8��tj P�L$<�%�Ë�$8  d�    Y_^[��]� ������U����j�h�Ad�    P��  SVW�  3�P��$�  d�    ��$<  �. ��$�  Ǆ$�      ���
 �L$LƄ$�  ��[���L$d��[���} u%�E����   ����$D  �$Q���҅��-  �]��u��$�  �E�؋�Bx���Ћ�����   �Ή|$$�Ѓ��D$8��  3���;��D$(%�D$,�D$0�D$4~W�L$,�<��3�;�Ƅ$�  |
;|$4�|$0��D$,�R|P���҅���  ����   ���ҋ��D$,� ����$�   �$Q��������$���D$,t�T$$����� ������L$$���T$��� ��$  �ʋ��������$R������D$����$,  �$P��������$$  Q��$  R��$�   P�����
 ����  ��t�H+�����$�{�
 �L$|Q���O�
 j ��$�   Ƅ$�  �S��� ����$�   �$R�����
 j��$�   ��R��� ����$�   �$P����
 ��$�   Q��������$�   R���������$�   P��$�   Qj j�6~
 �����  ��$�   R��$�   Pj j�~
 ������  ���U����Dz	��;�]�\$D�D$   �D$    �L$;L$$�N  �|$8�|?���|$}	�   �|$�D$3ۅ�����\$ݜ$�   �  �D$�D$,�L$��܌$�   ��$\  �������D��������$R������L$L�P�T$P�H�L$T�P�T$X�H�L$\�P�D$<P�L$PQ�M�T$h�7�
 ����   �D$D�D$<��������{p�M����$t  �$R�6�
 ��L$d�P�T$h�H�L$l�P�T$p�H�L$t�P�D$LP�L$h�T$|��o���]����At�D$<��;��\$D�\$�����
���D$    �D$�|$ ������L$|Ƅ$�  豟 �L$(Ƅ$�  ��;����$�  Ƅ$�   ���
 ��$<  Ǆ$�  �����u� �D$��$�  d�    Y_^[��]� �L$|Ƅ$�  �H� �L$(Ƅ$�  �w;����$�  Ƅ$�   ��
 ��$<  Ǆ$�  ������ 3���$�  d�    Y_^[��]� ��U����j�h�Ad�    P��(  SVW�  3�P��$8  d�    ���Ph�L$4Q���ҍL$4Ǆ$@      ��P������  �L$\��V���L$D��V����$�   ��V����$�   ��V����$,  �V����$  �V����$�   �V����$�   �V����$�   �V����$�   �V���E�}�T$|���\$t�D$3 ��   ��
{j �L$8�$O��� �]�L$4�����8  j�	O��� �]����Dz����   ���҅��1  ���L$4�  j �D$7��N��� jݜ$�   �L$8�N��� �\$t�6j �L$8�N��� �]������  j�L$8�N��� �]����A��  W��� �؍C������{  ���o�$��o�}�D$tW���S�L$dQ�����$�{�������   �D$|Wj�T$LR�����$�Z�����te�|$3 t0�D$D�L$H�T$L�D$\�D$P�L$`�L$T�T$d�T$X�D$h�L$l�T$p�E���$�D$LP��$�  Q�L$l��V�����y]������  �L$4��$@  �q� 2���$8  d�    Y_^[��]�8 �}�D$tW���S��$�   R�D$hP�����$������t��D$|Wj��$  Q�T$PR�����$�l�����t��|$3 t0�D$D�L$H�T$L�D$\�D$P�L$`�L$T�T$d�T$X�D$h�L$l�T$p�E���$�D$LP��$P  Q�L$l�V�����\����t7�E ���$��$  R��$�  P��$�   ��U�����k\������  �����$@  �L$4�`� 2���$8  d�    Y_^[��]�8 �}�D$tW���S��$�   Q�T$hR�����$������������D$|Wj��$�   P�L$PQ�����$��������n����|$3 t0�T$D�D$H�L$L�T$\�T$P�D$`�D$T�L$d�L$X�T$h�D$l�L$p�E���$�T$LR��$�  P�L$l��T�����[����������$�   Q��$�   �U���]0������  ������}�D$tW���S��$4  R��$�   P�L$lQ�����$�e�����������D$|Wj��$  R��$  P�L$TQ�����$�4������{����|$3 t0�T$D�D$H�L$L�T$\�T$P�D$`�D$T�L$d�L$X�T$h�D$l�L$p�E���$�T$LR��$h  P�L$l�T�����Z�����'����E ���$��$  Q��$�  R��$�   ��S�����[Z����������E(���$��$  ��$�  PQ��$<  �����}�D$tWj���$�   R��$�   P�L$lQ�����$�r�������   �D$|Wj��$�   R��$�   P�L$TQ�����$�A�����tU�|$3 u*�E���$�T$LR��$�  P�L$l�S�����Y����t$��$�   Q��$�   �(S���E0��������Au��Ǆ$@  ���������E8��$�   ��$�   ��(�\$ �ă����\$0���$�   �H��$�   �P��$�   �H��$�   �P��$�   �H��$�   �ĉ��$�   �H��$�   �P��$�   �H��$�   �P�Hu賝����@��u Ǆ$@  �����c���臜����@���4��������$@  �L$4��L$4Ǆ$@  ����蘗 ���$8  d�    Y_^[��]�8 ��j�j�l�kn�o �������̃�VW���L$�O���t$$���O���D$(j j V�D$P�����$�
���_��^��� U����j�hLBd�    P��  SVW�  3�P��$�  d�    ������}�\$<2ۃH����\$D����\$Lu9�GPj j �D$DP���$������u����\$<����\$D����\$L�G@=   �*  �L  ���F  �� �  ��$�   ���
 ��;����   ���$��$�   Pj ��Ǆ$�      �҄�tE�E��$�   ��$�   ���$�   �P��$�   �H��$�   �P��$�   �H�P��  3��D$T�$�D$X�D$\�D$`����   ��Ƅ$�  �҅���  ����   j �L$XQ���҅��|  �T$\���o  �|$X��E��O�H�O�H�O�H�O�H�O������H��   �r������ލLR��ۍύ��A0��`���T$<݁�   �T$D݁�   �T$L� ������@�X�@�X�Ax�T$<݁�   �T$D݁�   �T$L� ������@�X�@�X�A`�T$<�Ah�T$D�Ap�T$L� ������@�X�@�X�AH�T$<�AP�T$D�AX�T$L� ������@�X�@�X�D�����~>�R�ύ�    ����T$<�����A �T$D�A(�T$L� ������@�X�@�X��D$\�������� ������H�X�H�X��   �L$<�0V������   ��$$  �LL���L$|�CL���GPj j ��$�   R��$0  P�L$LQ�����$������tr�L$|�-S����������z\�ȍT$|��R�����$x  �$P�N����P��$@  Q�L$D�M����M��P�Q�P�Q�P�Q�P�Q�@�A���؍L$TƄ$�   �c�����$�   Ǆ$�  �����\�
 ��  ��$�   ��
 ��;����   ���$��$�   Pj ��Ǆ$�     �҄�t��L$|�1K���L$T�(K���D$TP��$�   Q��$�   ���
 ���t����T$<R��$�   �b���\$l�D$<P��$�   �qb���\$l�����D$|t�D$T�M���P�Q�P�Q�P�Q�P�@�Q�A�����=   tB�L$<�bT�����  �E�D$<��D$D�X�D$L�X���$�  d�    Y_^[��]� 3��D$T�$�D$X�D$\�D$`����   P�D$XP��Ǆ$�     �҅���   �D$X��u��P�V�H�N�P�V�H�N�P�D$<P�ΉV�ya���\$l�   9D$\�D$x�)  �D$X�   �L$<�Q���Ka���D$l������A�D$Xu0��\$l��L�N�T�V�L�N�T�V�L�N���؋L$x����;L$\�L$x|��   ��$T  R���������}��P�W�H�O�P�W�H�O�P�W����   �γ�҅�up�D$|P�������L$<Q���`���\$l�T$<R��$�   �|`���\$l����z8�D$|��$�   ��$�   ���$�   �O��$�   �W��$�   �G�O�W�D$X�|$` Ǆ$�  �����D$T�$t��tj P�L$\��$�Ë�$�  d�    Y_^[��]� �D$j ���\$�D$�$����� �����D$j ���\$�D$�$�W���� ���̋D$V��3�;���D�N�N�N~P��謻  ��� E^� j�hxBd�    PQVW�  3�P�D$d�    ��t$� E3��|$�&���9~�D$������Dt�F;�tWP����D�~�~�~�L$d�    Y_^����������U����j�h�Bd�    P���  SVW�  3�P��$�  d�    ��t$,��P43��ҋ���u�}���X���  �    �hY��  ��E���   �����$�҅���   �}���   �}  ��$  P�������P��$�   Q���M���P��$�   ��� �E���$W��$�   Ǆ$      ���
 ��u����$��$�   W���
 ��$�   Ǆ$   ������� ��  ����  ��Bx���Ћ؃��\$4��   ����   ���Ћ����|$x��   ��S�L$@�A�����Ǆ$      |
;\$H�\$D��D$@�R|P���҅���   ��Ph�L$dQ��������$�L$lƄ$  �>������$�   �$P����������$�L$l�>������$�   �$Q���������$�   �L����A����z?�L$dƄ$   ��� �L$<Ǆ$   �����")��3���$�  d�    Y_^[��]� ��~���|$(�D$(3��荌$�   ��|$8�\$|��D���L$L��D��9|$4�_�t  ���}  �D$@�D����\$�L$t���$�rO��3҅���;t$(�T$0�"  ���  �D$0�D$8Pj ܌$�   ��$�   Q���L$x�$�j=���L$8���$�{������������$�   R��$�   P��$�   �GF����L$L�P�T$P�H�L$T�P�T$X�H�L$\�P��$�   ��PQ�L$T�T$h�:F������$�   �$R�F����P��$  P�L$T��E����L$L�P�T$P�H�L$T�P�T$X�H�L$\�P�L$L�T$`��J����'����Az�   �3ۃ�;t$(�t$0������t$,��;|$4�������t��$�   P�L$P�C@���L$LQ��$�   R��$�   P��$P  �  �}��Ƅ$   t�    ��$D  �t$,�L$x�T	�T$(�D$(��$,  ��P��λ   ݜ$�   ��������̉�P�Q�P�Q�P�Q�P�@�Q�A��$�  ��N�����]����Au3�3��ۉ|$8��   ;|$4��   �D$@�D����\$�L$t���$�+M��3��ۉt$0��   ;t$(��   �D$0�L$8Qj ܌$�   ��$�   R���L$x�$�*;���L$8���$�;�����tX��$�   ��$�   ���ĉ��$�   �P��$�   �H��$�   �P��$�   �H��$�  �P�N�����]����Au3ۃ��ۉt$0�Q�������������$D  Ƅ$   �?� �L$dƄ$   �.� �|$H Ǆ$   �����D$<%t�D$@��tj P�L$D�%�Ë�$�  d�    Y_^[��]� �����V���H����D$t	V���������^� ��S�\$UVW���������GP��贴  �o3���~6�O�<� ���D$    t� ��ȋB�ЉD$�L$Q���� ��;�|�_^]�[� ������������V�t$��th8@���K�����t��^�3�^���������������̸8@�����������V�1��W|K�|$;�}C�Q��|<;�}8�A��|1;�}-�I��|&;�}";�t;�t;�t;�t;�t;�t
_�   ^� _3�^� �����̋D$VP��������u^� �F�@�W�|$�ύ@R���/B������   �F�@��ύ@R���B����tt�F�@�F�ύ@R����A����tX�F9FtW�@��ύ@R����A����t8�F�@�F�ύ@R���A����t�F�v�@�ύvR���A����u_2�^� _�^� ���������̉�8  ����������V��W�|$�FP���m� ��tA�N(Q���^� ��t2���   R����� ��t ��d  P���� ��t��  V���� _^� ���V�t$Wjj��h � @����m ����   S�GP���4� �؄���   �O Q���/� �؄�tz�W$R���� �؄�ti�G0P���� �؄�tX��0  Q���� �؄�tD�WR���� �؄�t3���  P���T~ �؄�t�O(Q����� �؄�t�W,R����� �؋��� ��u	[_��^� ��[_^� _��^� ���������̃�SVW���� �|$3��D$�D$�D$P�L$Qh � @��� �؄��Q  �|$�/  U�nU���N� �؄��  UhDE���������u#�`/�U �d/�E�h/�M�l/�U�D$P���� �؄���   �L$Q�_� ���T$R�ωF 轹 �؄���   �D$P詁 ���n0U�ωF$踺 �؄���   ���   Q��� ����؍�0  R��萺 �؄�t^�FP���O� �؄�tM���  Q���k� ���Ä�t6�|$|/�T$R���/� �؄�t�D$P�?� �F(����,V���n� ��]���� ��u_^��[��� _^��[��� ��������U������@����`   t/�E��P  �$�:5���\$0���E��@  �$�"5�������)�E��@  �$�5���\$0���E��P  �$��4���\$8���D$8��  �$�4���E����D$@��   �$�4���M���]�������̸    ��������������D$��������z�`E���\$�D$��XE���\$�D$�������������������D$��������D{C����������z�`E���\$�D$���\$�D$��XE���\$�D$���\$�D$����\$�D$�\$�D$�������̋A3�;A�����SVjh3ۋ�SV� ���V��V���V ��5�^�^(�^�^�^�^0�^��+�^�^8�^@��E�^D�VH�^`��^d�^P�F�F�F   �^X^[������������V���x����D$�^(3���N�V�N�D$�V��E������Au�A�3��وF����Az�   �3��V0�F�V8�N�VH�N@�VP�ND�^X^� ����D$���$�A2������t���\$����u�D$�\$�D$���$�2������t���D$��������Az���D$�D$������z
�ٸ   ���������Au����3���V3�W�|$8G����3�8N��+���  8G��3�8V��+���  8G��3�8N��+���  �F�O:�s_���^� v
_�   ^� ����\$�G�\$�F�$����������E  ����\$�G�\$�F�$����������  ����\$�G(�\$�F(�$����������   ����\$�G0�\$�F0�$����������   ����\$�G8�\$�F8�$�c���������   �N@�ɋG@3Ʌ�3�+���   �ND�ɋGD3Ʌ�3�+�u}��$���\$�GH�\$�FH�$�	�������uW����\$�GX�\$�FX�$���������u5����\$�GP�\$�FP�$���������u�v`�`;������;���_^� ������V��L$�FPjQ� 
 �VRjP� 
 �NQjP� 
 �VRjP� 
 �NQjP�} 
 �V(RjP�q 
 ��H�N0QjP�b 
 �V8RjP�V 
 �N@QjP�J 
 �VDRjP�> 
 �NHQjP�2 
 �VPRjP�& 
 ��H�NXQjP� 
 �V`RjP� 
 �NQjP��
 VjP��
 �VRjP��
 ��VjP��
 ��H^� �������V�t$Wj��j����� ����  �GSP����� �؄��2  �OQ����� �؄��  �WR����� �؄��  �GP���� �؄���   j ���� �؄���   �G�����$�)� �؄���   �G(�����$�� �؄���   �G0�����$��� �؄���   �G8�����$��� �؄�ty�O@Q���*� �؄�th�WDR���� �؄�tW�GH�����$�� �؄�tA�GP�����$�� �؄�t+�GX�����$�w� �؄�t� F�����$�^� �؋G`��|��~h�Eh�Ehx  h�E�G! ��3���t`P���� ��tV�GP���w� ��tG�Q���� ��t8�G�����$��� ��t$�WR���� ��t�GP���t� [_^� ��[_^� �����̃�SVW�������|$$�D$P�L$Q���D$    �D$    ��� �؄��  �|$�  �V�D$$P�ωT$(�Ű �|$$ �V�����ۈN�T$$t�D$$P��蠰 �؃|$$ �V���ۈN�T$$t�D$$P���{� �؃|$$ �V���ۈN�T$$t�D$$P���V� �؃|$$ ���ۈN��   �T$R���5� �؄���   �FP��谰 �؄���   �N(Q��蛰 �؄���   �V0R��膰 �؄���   �F8P���q� �؄�tt�N@Q���Я �؄�tc�VDR��迯 �؄�tR�FHP���>� �؄�tA�NPQ���-� �؄�t0�VXR���� �؄�t�D$P���
� �؄�t�N`Q���i� �؋F`��|��~#h�EhFh�  h�E�� ���F`    ��tj�|$|c�VR���"� �؄�tR�|$|KV���m� �؄�t=�FP��茯 �؄�t,�|$|%�NQ���$� �؄�t�|$|��V���,� ��_^��[��� ��������������̋��L$;�tB���A�X�Q�P�Q�P�A�X��0�A��X �A��X(��P0�Q�P4�Q�P8�I�H<� �VW�|$j��j���� ����   �P���;� ��ty�F�����$��� ��te�FP���� ��tV�NQ���	� ��tG�F�����$�� ��t3�F �����$�� ��t�F(�����$�m� ��t��0V����� _^� ��������̃���SUV��3��V�F�V��V �D$�V(�F�n�D$�F W�D$ �F(�^���L$ �T$�L$$�$���N0�D$4�L$8�Q;���|$0�D$P�L$Q���� ����   �|$��   �T$0R���D$4    �� ��ts�D$0P�׸ ��U�ω芭 ��tXS���� ��tL�L$Q���ެ ��t<�T$R���^� ��t,�D$ P���N� ��t�L$$Q���>� ��t�T$(R��议 _^][��� ����V��݆0  W���$�[(��������   ��ܞ0  ������   ݆8  ���$�,(��������   ��ܞ8  ������   ��@  ���*������   ��P  ����)������   ���=����$����up���y=����$����Az\����<����$����uH���Q=����$����Az4���(������$����{���(������$����z_�   ^�_3�^�����������̋��  ������������I��$����A{.����A��������u������(F������z�������� F����������V�t$��th�A���������t��^�3�^���������������̸�A�����������V�t$��th�B��軋����t��^�3�^���������������̸�B�����������V�t$��th�C���{�����t��^�3�^���������������̸�C����������̃���4F�A    �A�A���	 ������;������������̸   ����������̸   ����������̋A�I�T$PQhhGR詼 ��� ����������������̸   �����������V�t$Wh�GV���m� ������ h�GV�X� ��W���� h�&V�B� �GPh�GV�3� h�GV�(� ����螻 ��W���c� ���̻ ��腻 W���M� ��趻 ��读 _^� ����������j�h�Bd�    P��  �  3ĉ�$�  SV�  3�P��$�  d�    ��~����tA�L$�� �L$Ǆ$�      �D$,   腓 9F�L$��Ǆ$�  ������p �Ë�$�  d�    Y^[��$�  3��$� ���  ����V�t$Wjj��h � @����Z ��u_^� SW���6� �؄�t/�GP���5� �؄�t�OQ����� �؄�t�WR���� �؋���� ��u2ۊ�[_^� �����������̃�UVWh�   3���WV�*� ����V�D$�V@P�Vh�L$ݞ�   �n�|$�|$�|$Qh � @���� ��u	_^]��� �|$S�Ä���   V��蛩 �؄���   VhDE�6�������u"�`/��d/�F�h/�N�l/�V�FP���2� �؄�t>U���D� �؄�t0�|$|)�N�T$�L$R���� �؄�t�D$P�n ���F���g� ��u2ۊ�[_^]��� ����̸�D�����������VW�|$W���S ���   ���   ���   ���   ���   ���   ���   ���   W���   ���   �@m _��^� ����������T �����������V�t$Wj j��h � @���X ��u_3�^� ���   SP���� �؄�tL���   Q���
� �؄�t8���   R����� �؄�t$���   P���� �؄�t���   W���� �؋��� ��u2���[_^� �����̋L$h�G�½ �   � ���������̸�E�����������j�h8Cd�    P��SUVW�  3�P�D$(d�    ��l$�^Q ���   �E $H�   � A���D$�P��E�D$4    �|�����M�P�U�H�M�P�U� 0�E�0�M�0�U �0�E$�E(   �ƅ�    �ŋL$(d�    Y_^][�� ������������̸h   ����������́��   ���������V�t$Wj j��h � @����V ��u_3�^� Sj j h � @��2��J� ��t#V���   �*����ΈD$�/� ��t8\$t����� ��u2���[_^� ������������̃�SUV��W���   �   � A���|$,�D$P�L$Q3�h � @���E ƃ�    �t$ �t$(�4� ��u_^]3�[��� �|$�D$ uf�T$ R�D$P�ωt$ �t$(�t$,��� ��tE�|$ � @�D$, u9t$$|9t$ vW���B�����t�D$,����� ��t�|$, t�D$���� ��t�D$_^�E ]ƃ�    ��[��� ����������̋L$hdH�"� �   � ����������VW�|$��;~tfS3�;�~E9~~�~�N��PWQ����;ÉFt;�N;�~��+����R��SP��� ��[�~_^� �F;�t�SP�B�Љ^�^�^[_^� �������̋D$�L$�@��PQ�������� ����VW�|$��;~tjS3�;�~I9~~�~�N��PWQ����;ÉFt?�V;�~��+ʍI��Q�R��SP�O� ��[�~_^� �F;�t�SP�B�Љ^�^�^[_^� ���̋D$�L$PQ�Q������ �����������S�\$��V��~SU�l$��|IW�|$��|?;�t;�F�+;�1;�-�N�;�~�;�}��P���6����F�(SR�P�&� ��_]^[� �����������̋D$�T$��    QR������� ���̋D$�L$��PQ������� ��������VW�|$��;~tlS3�;�~K9~~�~�N��PWQ����;ÉFtA�V;�~��+ʍI���Q�R��SP��� ��[�~_^� �F;�t�SP�B�Љ^�^�^[_^� ��SW�|$����~dU�l$��|ZV�t$��|P;�tL�C�/;�B;�>�K�>;�~�;�}��P���6����C����R�Lm ��R�v��R��� ��^]_[� �����������S�\$��U��~[W�|$��|QV�t$��|G;�tC�E�;�9;�5�M�;�~�;�}��P���V]���E����S����WV�n� ��^_][� ���̋Q2���t(�I��~!V�t$��t��~Vh�   QR��d ���^� �����������̋Q2���t(�I��~!V�t$��t��~Vh�   QR�d ���^� �����������̋D$�L$i��   PQ������� �����V���������h  �X  ���   �p  �  N$�J�NDN4N�I�Q��x  ����H  �  ^������������V��F�N�@Q�L$��PQ�$
 �V�N R��QP�
 �N,�v0�v�Q�RP��

 ��$^� ������̃��  3ĉD$�D$=   SUV�t$(W��}�   �3�=   �Í\S��� � �˃���   ��tO���
  3�9\$(��   3����   �G�Pj��貮 ����;\$(|�_^][�L$3��Q� ��� 3�9\$(��   3�I ����   �G�(�f�L$�Pf�T$�Hf�L$�P�D$Pj��f�T$"衬 ����;\$(|�_^][�L$3���� ��� 3�9\$(~K3퍛    ��t?�G�(ňL$�P�T$�H�L$�P�D$Pj�ΈT$詫 ����;\$(|��L$_^][3��x� ��� �������̃��  3ĉD$SU�l$,VW�|$0��3�9{$�t$}	W�K�0Z���D$P��脜 �L$����   ��tA����   3�;���   �t$����   �CD$��Pj�2� �D$��;�|��   3�����   �t$�I ����   �L$Qj���Z� �KL$�T$�D$��T$�Q�T$ �Q�T$"��;��Q|��N3���~H�t$��t@�D$Pj��蚠 �KL$�T$�D$��T$�Q�T$�Q�T$��;��Q|���|;s$�s �L$$_^][3��� ��� ������̃�SV��L$W�z �|$�ȋF;��L$�~_^2�[��� ����  3�;F0U��3ۃ�#�;��   ����3҃�#�;�l  �\$��#׉T$ 3�;�  ��#׃��T$ue�FPP�jP�l �F,PP�Lm jQ�l ���   PP�jR��k ��h  PP�D$X� jQ��k ��  �T$P��@PPjR��k ���F�L$$P���P�.�
 �؄�tz�F,�Lm ��PQ�L$,��
 �؄�t^���   �T$�L$$P��    P���
 �؄�t<��h  �L$ ��PQ�L$,���
 �؄�t��  �T$�L$$P��    P��
 �؃|$ui�FPP�jQ�k �F,PP�Tm jR�k ���   PP�D$<� jQ��j ��h  �T$PPP�jP��j ��  �L$P��@VVjQ��j ��]_^��[��� ��V��~ �lIt%�F��tj P�xI�F    �F    �F    ^�����������VW�|$��;�t>�G��_�F    ��^� 9F}P�����N��t�G�F��P�GPQ�9� ��_��^� ���������������S�\$��V��~[U�l$��|QW�|$��|G;�tC�F�+;�9;�5�N�;�~�;�}��P�������F��    R��Q��R�.� ��_]^[� ����VW�|$��;�tA�G��_�F    ��^� 9F}P�4����N��t�G�F�W���PRQ�f� ��_��^� ������������QU�l$V��W���w �|$���D$��  S�D$P���D$     ��
 �؄�t`�D$��tX���;�u/�NW�F����F�T$RP�D$$P���A�
 �؄�t)W�N��T���h�Jh�Jh�  h�E� ��2ۄ��D$    tr�L$Q���*�
 �؄�t`�D$��tX���;�u/�N(W������F,�T$�L$QPR�����
 �؄�t)W�N(�tT���h\Jh�Jh�  h�E� ��2ۄ��D$    t{�D$P����
 �؄�ti�D$��ta��    ;�u8���   W�������   �T$RP�D$$P���?�
 �؄�t,W���   ��S���hJh�Jh�  h�E� ��2ۄ��D$    ty�L$Q���%�
 �؄�tg�D$��t_����;�u8��d  W�������h  �T$�L$QPR����
 �؄�t,W��d  �hS���h�Ih�Jh�  h�E�} ��2ۄ��D$    t{�D$P����
 �؄�ti�D$��ta��    ;�u8��  W苌  ��  �T$RP�D$$P���3�
 �؄�t,W��  ��R���h�Ih�Jh�  h�E�� ��2ۃ|$uu�FPP�F�@jQ�wf �F,PP�F0�@jR�df ���   PP���   �jP�Lf ��h  ��l  PP�jQ�4f ��  ��  ��@PP�vjR�f ����[_^]Y� �����������V��L$��|-�F;�}&+���P�APQ��������F��N�V3��ʉ�A^� ����SW�|$����~bU�l$��|XV�t$��|N;�tJ�C�/;�@;�<�K�>;�~�;�}��P��������C���R�Lm ��R�v��R��� ��^]_[� �������������V��L$��|3�F;�},+���P�APQ���\����F��N�V3��I����A�A^� ��������������V��~ ��Ht%�F��tj P��H�F    �F    �F    ^�����������VW�|$��;�t;�G��_�F    ��^� 9F}P�����N��t�GP�F�GPQ�|� ��_��^� ��V��L$��|(�F;�}!+���P�APQ���<����F��F�N�� ^� ���������V��~ ��Ht%�F��tj P��H�F    �F    �F    ^�����������V��~ ��Ht%�F��tj P��H�F    �F    �F    ^�����������V��~ ��Ht%�F��tj P� I�F    �F    �F    ^�����������V��~ �It%�F��tj P�I�F    �F    �F    ^�����������VW�|$��;�tB�G��_�F    ��^� 9F}P�} �N��t�G�F�W����PRQ��� ��_��^� �����������V��~ �It%�F��tj P�(I�F    �F    �F    ^�����������V��L$��|<�F;�}5+���P�APQ�������F��N�V3��I�ʉ�A�A�A�A�A^� �����V��~ �0It%�F��tj P�<I�F    �F    �F    ^�����������VW�|$��;�t>�G��_�F    ��^� 9F}P�N���N��t�G�F��P�GPQ�� ��_��^� ���������������V��L$��|3�F;�},+���P�APQ�������F��F3���F��H�H�H^� ��������������V��~ �XIt%�F��tj P�dI�F    �F    �F    ^����������̋A��~9A0u��2���������������̋A��~9��   u��2������������̋A��~9�  u��2�������������SVW���  �   ���7��t�N0�"Z V�<������    ����u�_^[��������U������SVW�y��~o9y0uj�I,j ��,���L$���1����~F��L$�\$�F�\$�F�\$ �p����u2��D$���^����D$�����^��D$ �^�u���_^[��]�_^2�[��]������W���G��~*9G0u%��~!SV3��؍�$    �O,��������u�^[_�����������V���������^����̋���������V3��V0�F�V8�F�VH�FD�VP��^X�F��E�F�^�F@   �5�F   �^(�����������������̋��i������V3��V0�F�V8�F�VH�FD�^P�� K�F�^�F�5�F@   �^(�F   ��E���^X����������V�������F(���\$����$�$�n����F   ^������j�hkCd�    PQVW�  3�P�D$d�    ��t$�~0���	�����V3��V���V ���V(�D$(�T$��$�F�F�����ƋL$d�    Y_^���������������U����j�h�Cd�    P��hSVW�  3�P�D$xd�    ��}3�;�~9Et��\$7��D$7������V�N0�V��V �F�V(�F�T$�$�N������  �L$<�M� W�L$@Ǆ$�       �H� �؋E�P����T$8wE�$�����E��������At���K�^�$���E��������At���K�^��D$7 ����   �M����wa�$�(��A�	�U�A���$���F����A��������Az������(F������z���������� F������������������^����u�F���1�V��t�V0����{�V8����Au�V8��V8�V0�ӃF�T$8�����E����F��u2��   PSj�U �N���+����Ë�� ����  ��V�L$8yJ���Bu�@���$�������^���3���~�Ã�;��F �^ |��D$83����F ���V ~�Ã�;������F(�^(|��؊\$7�~(�^(�L$<Ǆ$�   �����2� �ËL$xd�    Y_^[��]� �I @�_�_�_����������������V��~ ��It%�F��tj P��I�F    �F    �F    �D$t	V�ߟ������^� ������V��~ ��Jt%�F��tj P��J�F    �F    �F    �D$t	V菟������^� ������V��~ ��Ht%�F��tj P��H�F    �F    �F    �D$t	V�?�������^� ������V��~ ��Ht%�F��tj P��H�F    �F    �F    �D$t	V��������^� ������V��~ ��Ht%�F��tj P��H�F    �F    �F    �D$t	V蟞������^� ������V��~ ��Ht%�F��tj P� I�F    �F    �F    �D$t	V�O�������^� ������V��~ �It%�F��tj P�I�F    �F    �F    �D$t	V���������^� ������V��~ �It%�F��tj P�(I�F    �F    �F    �D$t	V话������^� ������V��~ �0It%�F��tj P�<I�F    �F    �F    �D$t	V�_�������^� ������V��~ �XIt%�F��tj P�dI�F    �F    �F    �D$t	V��������^� ������U��������  ݁0  ��  ݁8  Sݙ0  ��   Vݙ8  ��  W��  ��  ��$  ��  ��(  ��  ��,  ��   ��$  ��(  �t$��  ��,  �|$3�����  ��  �D$�T$|Q�V������A(�<�    ��    �@؃�@���@��X��X��@��@��X��X��@��@��X��X��@��@��X��X�u�;�}�����+�� �����@��X��X�u�L$�P _^�[��]�������U����j�h�Cd�    P��   SUVW�  3�P��$�   d�    ��F��~���   ;�l$Ht2���$�   d�    Y_^][��]�������~\ �~H��uW��������u��������t�����  ����  ��@  �������P  �͊����:��À�`   t����h@h`�jj�D$tP�q  ��W�G�L$d�O�T$h�U �L$p�M�D$l�E�T$t�U�L$|�L$dǄ$�       �D$x��$�   �~���L$t�u��3�9l$H��   ���   ��<�    �L$T�T8j �L$X�T$\�b��� ���L$l�$�� ���\$Lj�L$X�B��� ���L$|�$� ����u���D$L���\$L����L$l�$�@ ���\$\�D$L���L$|�$�) ���\$L�D$L���   ���\$��D$d�\$T�D$T�$������;l$H�8���h@jj�D$pPǄ$�   ������� ��   3Ƀ���   �}����   ��    ���\$H���@��D$H�X���   �D�D�\$H���@��D$H�X���   �D��D��\$H�@��D$H�X���   ��;��\$H�@��D$H�X�y���;�}(��I ���   �ʍ��\$H��;��@��D$H�X|ݰ��$�   d�    Y_^][��]�����U����j�hDd�    P��hSVW�  3�P�D$xd�    ��}���  �F����  9��   ��  ������~\ �^H�D$+uS��������u��������t��|$+ ���   �\$,��   ����   ��`   t	�   +ǋ��O���1�D1ΉT$4�Q�D$8�A�T$<�D$@3ۉ�$�   ����9\$,~S���   ��W�L$4����� ���L$<�$�'���������L$<�$�������t	�T$0�Z��D$0���;\$,|��L$4Ǆ$�   �����TL ��L$xd�    Y_^[��]� ��3҃���   ������   ��    ���t
�@���X�� ��������   �Dt
�@���X�� ������   �����D�t
�@���X�� ������   ���t
�@���X�� �����;��w����\$,;�}$�����   ��t
�@���X�� �����;�|��ذ�L$xd�    Y_^[��]� 2��L$xd�    Y_^[��]� ��������VW�|$�����  �F���  9�  �  �GS���0U���V�����t���������  3�����   �]���3Ƀ���    �T$�d$ ��  ���t
�@���X�� �������  �Dt
�@���X�� �������  �Q0�D�t
�@���X�� �����  �t
�@���X�� �����@��u��D$;�}-����+�Ջ�  ���t
�@���X�� �������u�][_�^� _2�^� ������������j�hIDd�    PQSVW�  3�P�D$d�    ��h���D$    �L$(h���D$$    �WI ����D$    �D$   ��   �D$(����   ;G,��   ��G(�ȋ��|y�W;�}r�I��|k;�}g�W�����ʃx ~T�@��tM�y ~G�I��t@� ���1�K|5;�}1��|-;�})�K�\$$�@��R���u����P�v��P�K�a���D$$�L$d�    Y_^[��� ��������j�h{Dd�    PQV�  3�P�D$d�    j�ב�������t$���D$    t0�����	 ����F�F�4F�F    �ƋL$d�    Y^���3��L$d�    Y^������������������j�h�Dd�    PQVW�  3�P�D$d�    ��j�D��������t$���D$    t$���h�	 �4F�F    �F�����F�����3����D$����t;�tW���q�	 �G�F�O�N�W�V�ƋL$d�    Y_^��������������VW�|$��tKh�A���]����t;�t$��t3h�A���]����t#;�tW����	 �G�F�O�N�W�V_�^�_2�^�������j�h�Dd�    PQV�  3�P�D$d�    j�7��������t$���D$    t.���[�	 ��F�F    �F�����ƋL$d�    Y^���3��L$d�    Y^����j�hEd�    PQVW�  3�P�D$d�    ��j贏�������t$���D$    t���ث	 ��F�F    �F�����3����D$����t;�tW����	 �G�F�O�N�ƋL$d�    Y_^�����������VW�|$��tEh�B���\����t5�t$��t-h�B���\����t;�tW��肫	 �G�F�O�N_�^�_2�^�������������j�h;Ed�    PQV�  3�P�D$d�    j跎�������t$���D$    t.���۪	 �G�F    �F�����ƋL$d�    Y^���3��L$d�    Y^����j�hkEd�    PQVW�  3�P�D$d�    ��j�4��������t$���D$    t���X�	 �G�F    �F�����3����D$����t;�tW���h�	 �G�F�O�N�ƋL$d�    Y_^�����������VW�|$��tEh�C���Z����t5�t$��t-h�C���Z����t;�tW����	 �G�F�O�N_�^�_2�^�������������V�����4F�F    �F�F��	 �D$t	V�5�������^� �����������̋A��u�D$��thLP趋 ��3�� W�y���t*��|;x|C�L$��t�@PWh�KQ脋 ��3�_� �y�u�D$��th�KP�b� ��3�_� V�q�����   ��8  ��u�D$��tVh�KP�.� ��^3�_� ��|Q;q,}L���ti����A3ɋP��~�@��98t
����;�|�;�|A�D$��t2VWhXKP�ي ��^3�_� �D$��t�IQVh$KP跊 ��^3�_� ^�   _� ��̡��V�t$�����V����F����V����F����V�Q��tE�A���u#�A��|6;�T  }.���P  �x ~�@� ��|;B}�R�@��P��������^� �������V����F�F    �F������	 �D$t	V�7�������^� �������������̋Q��u�D$��tHhLP趉 ��3�� �A��|;�d  }�   � �L$��t��d  RPh,LQ�|� ��3�� ����V���G�F    �F�����D�	 �D$t	V藌������^� �������������̋Q��u�D$��tBhLP�� ��3�� �A��|;B }�   � �L$��t�R RPh\LQ�� ��3�� ���������̃�dSU�ًSV2���W��   �K����   ;J ��   h���P��Hjj�D$ P�T$ ���I��3��|$�D� ��|^;D$}X�S�@�B��Q�������������|ӋD$|�L$x3�9�$�   ��RPQ�T$ Rjjj j�6N �� _^]��[��d� _^]3�[��d� ����������VW�|$j���j ���m�
 �F��|�v��t;F}<Pj����
 ��_^� �F��|$�v��t;F}��T  ��t;�}
Pj��训
 ��_^� �������VW�|$j���j �����
 �F��|�v��t��d  ��t;�}
Pj���g�
 ��_^� VW�|$j���j ��轫
 �F��|�v��t;F }
Pj���0�
 ��_^� ���������SV��W�~������h�   3�SV�� ������V@_�Vh��ݞ�   ���   ���   ���   ǆ�   �H���   ^[���������VW�|$��t5h�D����T����t%�t$��th�D����T����tW�������_�^�_2�^�������������j�h�Ed�    PQSVW�  3�P�D$d�    ���|$��L3�9��   ���   �\$��$t�F;�tSP����$�^�^�^���D$�����}  �L$d�    Y_^[������������̋��   V�4@�����! �^��������V��L$���   PjQ��	 ���   RjP�{�	 ���   QjP�l�	 ���   RjP�]�	 ���   ���   �v��Q�RP�@�	 ��<^� ���������U������ VW���L$�����D$P��D�P��P���CQ������th�D���AS����u2�_^��]ËW;��   u�ҋ���   tJ����\$�A�\$�A�\$�D$�������Dz��D$�G������Dz��D$�G������Dz���u�_�^��]�����������̃�V�D$��P��D�P��P���P������th�D���R����u3�3�����^�����������������̋D$�H�@�@�Q�Rj ��	 ����̃�VW�D$��P��D�O��P���"P������t8h�D��� R����t(�N���   �V�v�v�R�Pj ��	 �����   _^����������������̃�V�D$��P��D�+O��P���O������t?h�D���Q����t/���   ���@����   ���   �R�Pj �7�	 �����   ^�����������̃�VW�D$��P��D�N��P���BO������th�D���@Q����u_�^��Ë��   ;Nu,�V�v�v�R�Pj ���	 ��9��   u_�   ^���_3�^�������̃�V�D$��P��D�;N��P����N������th�D����P����u�^��Ë��   ;��   u3���   ���   �@��R�Pj �:�	 ��9��   u
�   ^���3�^�����������������j�h�Ed�    PQ�  3�P�D$d�    h   �E������D$���D$    t�������L$d�    Y���3��L$d�    Y������������j�h�Ed�    PQSVW�  3�P�D$d�    ��h   �Ђ�����D$���D$    t���&������3ۅ��D$����tV��� �Ƹ   ���   �   �ËL$d�    Y_^[�������V�t$��WtHh�E���JO����t8�|$��t0h�E���2O����t V���& �Ƹ   �Ǹ   �   �_�^�_2�^����������j�h+Fd�    P��VW�  3�P�D$d�    �|$,��u3��L$d�    Y_^��ÍD$P��E�L��P���L������th�E���N����u?3��|$0 t6h   菁�����D$,���t$$t	��������3�P���D$(��������S���ƋL$d�    Y_^������������������V���$H�r �D$t	V�%�������^� ������������jQ���������u2�� V�t$W���   �   ��󥋈�   ��_�ƀ�    ^t��t
ǀ�      �� ������������V��~ t&�F��t�j P�B���F    �F    �F    ^����������������j�haFd�    PQ�  3�P�D$d�    �L$�L$���D$    t������L$d�    Y��� ����V��~ ��Ht%�F��tj P��H�F    �F    �F    ^�����������V��~ ��Jt%�F��tj P��J�F    �F    �F    ^�����������V��~ ��It%�F��tj P��I�F    �F    �F    ^����������̃�SUV�t$Wj��j����� �o �؄ۋG�D$�l$��   P���| �؄���   U���| �؄���   ��@  P���.� �؄���   ��P  Q���� �؄�t|��  R���� �؄�th��   P���� �؄�tT��0  Qj���{ �؄�t>���  Rj���r{ �؄�t(���  Pj���\{ �؄�t���  Qj���F{ �����  ����� t��t	��u3��
�   ������t
Q���!{ �؃��   �D$ ��tH�T$ R����x �؄�t6�|$  t/j h � @��� �؄�t���  V趶���Ί�轥 ��u2ۄ��D$    ��   ���  ��|$}X�}  ���D$ �D$ P�dx �|$  ��t,j h � @��� �؄�t�M V�����Ί��U� ��u2ۃD$����u��+��t'�L$�T$VQR��������؄�t�D$VP���������3�8�`  ������   P���z �؄���   �GHP����{ �؄���   �L$��~o��  3�;��΃�#Ћ��	H ���D$ u��  PP�D- jP��9 ����  ����PQ���e�
 �|$ ��u��  PP�T- jR��9 ����tJV�OH������؄�t;���  P���#w �؄�t&���  Q���w �؄�t���  R����v ��_^]��[��� ������������ّ�  ّ�  ّ�  �hEّ�  ّ�  ّ�  ّ�  ّ�  ّ�  ّ�  ٙ�  ّ�  ّ�  ّ�  ّ�  ٙ�  �S������SV��W�s3�9~t�F;�t�WP�B���Љ~�~�~9{ �st�F;�t�WP�B���Љ~�~�~9{0�s$t�F;�t�WP�B���Љ~�~�~9{@�s4t�F;�t�WP�B���Љ~�~�~�sD;�t��    �Ƌ6P�f�����;�u�KH����{Dt�{H_^[��������������j�h�Fd�    PQVW�  3�P�D$d�    �L$3�9y�q�|$t�F;�t�WP�B���Љ~�~�~9~�D$�����It�F;�tWP���(I�~�~�~�L$d�    Y_^���̃�VW�|$$��F�N�VPQRh�LW��x ���D$P���/����L$�&�����t6���;x h�LW�x ���L$Q���{ h�&W�x �����Lx _^��� ���̃�S�D$P2�������L$�������t3�T$$�D$ 3�9L$(��QRP�L$Qjjj j�M> �� ��[��� ��[��� ������j�h�Fd�    P��0SUVW�  3�P�D$Dd�    ��3ۉ\$�t$Th��h���Ή\$T�/ �G;É\$L�D$   �6  �O;��+  ��8  ;��  ;A,�  ��A(���  �L$��	 ����D$4F�\$$�M �G�T$,�L$(R�L$�D$P   �D$$�������P�V�H�N�P�V�H�N�P�ΉV������tw�E�L$,Q�L$�D$,�s�����V�P�N�Q�P�Q�P�Q�P�Q�@�A�H�����u3��������V����F����N����V����F�L$�D$L �D$4F�D$     �\$$�\$(�{�	 �ƋL$Dd�    Y_^][��<� ���j�h�Fd�    P��  �  3ĉ�$�  SUVW�  3�P��$�  d�    ��L$�M �=`/�d/�-h/�l/h�   j VǄ$�      �D$@   �|$(�\$,�l$0�D$4�s� ��L$4�V�>�V@�^�Vh�nݞ�   �N���L$�F   ��M �L$�FǄ$�  �����+ ��$�  d�    Y_^][��$�  3��b� ���  ��j�hFGd�    P��V�  3�P�D$d�    ��t$� 3����   �D$$��L���   ���   ���   ���   �r( �D$P��D�D$(�@����N�P�V�H�N�P�V� 0�F�0�N�0�V �0�F$�F(   �ƋL$d�    Y^�� ������������V���8����D$t	V��w������^� �̃�SUV���   W3��8�D$���   ���   ���   ���   �;�} �89~�D$t�F;�t�WP�B���Љ~�~�~�L$Q�T$�|$�|$�|$(Rh � @��趫 ��u_^]3�[��� S���.a �؄�t<U��� a �؄�t.�D$P���a �؄�t�L$Q����` �؄�t
V���~j �؋��e� ��u2�_^]��[��� ��V�񋆼   9��   t h�Mh�Mhj$  h�E�V� ��3�^�;��   t h�Mh�Mhp$  h�E�.� ��3�^Ë��   P���   �@���Qj �	�	 ��9��   t h�Mh�Mhv$  h�E��� ��3�^�W��� ����th8@���A����u!h`Mh�Mh}$  h�E�� ��_3�^Ë��   ;Wt!h@Mh�Mh�$  h�E�{� ��_3�^Ã�W�J�����9��   t!hMh�Mh�$  h�E�F� ��_3�^�_�   ^���������U�l$W�������$�q������   ���   SV���   P�F�@���Qj ���	 ��U�΋��� �V�v�v��R�Pj ���	 ��;��   ^[u���   ;��   u���   _�   ]� 3҅����   _�   ]� �������U������SUVW��D$P��D�=��P���=��������   h�D���?������   ���   9}�]}W���&�����|;{�{���E���   t�������A�����X��A��X�u㋆�   ���   ���   �C�K�@�Q�Rj ���	 ���   ���   P���   �@���Qj ��	 �����   _^][��]����U������(SUVW���D$(P��D�|$�<��P���<���؅��B  h�D���>�����.  �o;��   ���   �D$9n}U���'�����|;n�n�|$ ���   �ts�L$��������   ����\$�F�\$ �F�\$$�D$�������Dz �D$ �G������Dz�D$$�G������D{���G�^�G�^������u��%��t!�d$ �������G�����^��G��^�u�D$�H���   �P���   �H�@�@�Q�Rj �G�	 ���   ���   P���   �@���Qj �#�	 �����   _^][��]��̃�SV��F�V;�W�|$ ��   ������   v��|� � ;�}�ȍ����   ~� �N��to��+���xf;�}b�L$�J���9^��G�O�T$�W�D$�L$�T$}S��蒕���F�L$��F_��T$�P�L$�H�T$�P�F^[��� ;�}S���U����F���F��W�P�O�H�W_�P�F^[��� ��������̃�S�\$V��F�V;�W��   ��    ��   v��|�  ;�}�ȍ<����   ~�< �N��tR��+���xI;�}E�L$�H���9~��C�T$�D$}W�������N�F�T$�ȋT$_�T��F^[��� ;�}W���������N�F�ȋS_�T��F^[��� �VW�|$����~V�|$ tO�FSU�n�8;�~詽��;�}��;�}P�������F�T$����Q�NR�@��R薲 ��~][_^� ��������̃�SUV��F�n;�W�|$ ��   �@�Ɂ�   v��|���� ;�}�ȍ����   ~� �F��tr��+ȸ���*���������x\;�}X�L$�����9^��G�O�T$�D$�L$}S���9����F�L$�@�F����T$�P�L$_�H�F^][��� ;�}S��������F��@�F����W�P�O_�H�F^][��� �����V��F�V;�u;������   v��|� � ;�}�������   ��;�}P���x���F��F3ɉ�H�H�H�N����F���N^���������������̃�$�D$,� S�\$V�@���\$�L$�@�\$$�(����D$$���\$@�L$�D$@���\$�D$(�\$@�D$@�\$�D$ �\$@�D$@�$�����D$0���N0|D;�}'�N,�T$�@����L$�H�T$�P^��[��$� u�D$P�N(�����^��[��$� ^2�[��$� ���D$V�\$���D$���\$�L$�D$�\$�D$�$�����L$���   2���|3;�}���   �D$�΋T$�T��^� u�D$P���   �����^� �����������j�h�Gd�    PQSVW�  3�P�D$d�    ���|$�D$   �����w43�9^�D$�It�F;�tSP���I�^�^�^9_0�w$�D$��Ht�F;�tSP��� I�^�^�^9_ �w�\$��Ht�F;�tSP����H�^�^�^9_�w�D$������$t�F;�tSP����$�^�^�^�L$d�    Y_^[�����������������j�h�Gd�    P��0VW�  3�P�D$<d�    ���G�O�t$LPQh�MV��h ���T$R�������L$�D$D    ������tP���'h h�LV�h ���D$P���mk h�MV�h ���L$$Q���Sk h�&V�hh �����h �L$�D$D�����}  �L$<d�    Y_^��<� ���������j�h�Gd�    P��0SV�  3�P�D$<d�    �D$P3�������L$�\$D�R�����t7�L$$�E�����t*�T$P�D$L3�9\$T��QRP�L$QjjSj��- �� �؍L$���D$D������ �ƋL$<d�    Y^[��<� �������������j�h+Hd�    PQ�  3�P�D$d�    h�   �h�����D$���D$    t��������L$d�    Y���3��L$d�    Y������������j�h[Hd�    PQVW�  3�P�D$d�    ��h�   �1h�����D$���D$    t���W������3����D$����tW���-����ƋL$d�    Y_^������������j�h�Hd�    P��VW�  3�P�D$ d�    �D$P��D��1���|$0P���2��3�;�t$h�D���~4����t3��L$ d�    Y_^�� �h�   �lg�����D$;Ɖt$(t	��������V���D$,�����9���ƋL$ d�    Y_^�� Ã�VW�D$��P��D�j1��P����1������th�D����3����uW�������ϋ������_���   ^��Ë��   ;��   u)���   ���   �@��R�Pj �R�	 ��9��   t3���   ;Ou(�G�W�@�R�Pj �&�	 ��9��   u������_���   ^�����������U������4�ESVW���W �O�؀�������\$�D$�T$$�L$}5��th�PP��d ����t2���_^[��]� 賿 ��_^[��]� ��}��t�h�P�ċw0��~;�t��t�QVhPPP�{d ��묋��   ��~;�t��t�QRhPP�Wd ��눋�  ��~!;�t���r���QRh�OP�/d ���]�������   ;���   ���D$     ��   3���I �G,�4j�������\$(j�������L$(j ���\$4�����j �\$,��������L$(j���D$4�\$,�����j�\$4��������L$0�D$(�\$(�D$(��O�����  ��O����A�  �D$ �؃���;D$�D$ �X���3����  �C���$�b��������  ����$�J���������   ������|čT$03�R��D�t$$�.��P���'/������  h�D���#1������  ���$������D$t��������p�t$ �������ϊ��n�������   �|$ ��   ����   ����   �D$��tqh�OP�xb ��8\$�����t$��t0�Ϡ �\$(�D$(�L$ ���$QhHOV�Ab ���|$ �l����|$ ���`����D$��thOP�b ���|$ �@����D$��t�h�NP��a ���|$ � ����D$��t�h�NP��a ���|$ � �������   3�9t$$~,3ۍ�    �D$ �O�T$P�R������t����;t$$|ܸ   _^[��]� �\$��t=�D$����OP脑����VuhTNS�Ta ���|$ ����hNS�<a ���|$ �g����\$$3���~�����L$Q���4�����t����;�|�_^�   [��]� �D$��t�VhTNP��` ���|$ �����������U������tSVW���G �w�L$P�D$<�t$8�;����L$h�2�����~;�L$@Q��D�/,��P���,����t h�D���.����t���,������D$7u�D$7 �W �G�uRPh�SV�H` ���|$7 �tEu�lEPh�SV�(` �G����~
9G0�tEt�lEPh�SV�` �G ����~
9G@�tEt�lEPhpSV��_ �G����~9�  �tEt�lEPhXSV�_ �G����~9��   �tEt�lEPh@SV�_ �G����~9�l  �tEt�lEPh(SV�f_ �G����~9�  �tEt�lEPhSV�>_ hSV�3_ �����^ V��x  蝢������^ ��`   �tEu�lEPh�RV��^ ����P  j���U������$j ���F������$��@  j���1������$j ���"������$h�RV�^ ��(��   j����������$j ����������$��  j����������$j ����������$h�RV�K^ ݇0  ���\$݇0  �$h�RV�*^ h�RV�^ �� ���] V�OH茡������] ���~] �OQhlRV��] �����e] �|$7 �D$@    t��������P�T$@�D$83ۅ���   ��u��~hdRV�] �\$@������   �O�[��R�L$T�����|$@ te�L$@�[�����T$h��0�@ݔ$�   �@ݔ$�   �\$(�\$ �\$݄$�   �\$݄$�   �\$݄$�   �$Sh,RV�] ��<�)�D$`���\$�D$p�\$�D$h�$ShRV��\ ��$�D$8��;��%������\ �O����   �G0;���   Ph�QV�\ �����,\ 3�9\$8~l�D$8��u��~hdRV�\ �\$@������<�G,�[��Q�L$T������D$`���\$�D$p�\$�D$h�$Sh�QV�F\ ��$�D$8��;�|�����[ �O����   ���   ;���   Ph�QV�\ �����[ 3�9\$8~t�D$8��    ��u��~hdRV��[ �\$@������>���   �؋D��T$@�D$@�T$P���D$T�D$T�T$h�\$�$Sh�QV�[ ���D$8��;�|����?[ �O����   ��  ;�u}Ph�QV�^[ ������Z 3�9\$8~X��u�|$8~hdRV�5[ �\$@������,��  �������@���\$�$ShlQV� [ ����;\$8|����Z �W Rh\QV��Z �����TZ 3�9\$<��   �D$<�d$ ��u��~hdRV�Z �\$D������V�O�����T�;Q�Ou�T��HR�QRSh@QV�oZ ���!�T��HR�P� QRPSh$QV�LZ ���D$<��;��z�������Y �O ����   �G@;���   PhQV�Z �����Y 3�9\$<~h��u�|$<~hdRV��Y �\$D������<�W<�[��P�L$T�Y����D$`���\$�D$p�\$�D$h�$Sh�PV�Y ��$��;\$<|����PY ���IY _^[��]� U����j�h�Hd�    P���   SVW�  3�P��$�   d�    ��N �V3����T$�0  ���'  �L$� ن�  ن�  ���  ���  ��Ǆ$       �����  ���n�������   ���/�������   ��������@j �L$hQ�T$TRP�D$(jPj j�� ���� ����   �D$L���$賍����D$\�$襍���_�D$d�$薍���_�D$l�$�Ǎ����D$t�$蹍���[�D$|�$認�����[��������tG�N�T$jSWQjRj j�# �� �*�Fj SWP�D$(jPj j�d# ���� ���D$��   ��L$�\$ن�  �\$$ن�  �\$,��\$4ن�  �\$<ن�  �\$D���������D$��   �} �u�}tSV��$�   �����W�L$P������L$|Q�T$PR��$�   �= P�L$ Ƅ$  �� ��$�   Ƅ$    �w �D$��D$$�_�D$,�_�D$4��D$<�^�D$D�^�L$Ǆ$   �����; �D$��$�   d�    Y_^[��]� ���������������SV3�8\$W��tO���  ;�t���2���W�Z�������  ��8  ���F������  ;�tP��Y�������  ���v����2��8  ��_�_�_�_�_ �_�_,�_0�_(�_<�_@�_8�_D�_H���{������  ���  �7��4  ���  ���  ���  ���  ���  ���  ���  _���  ^[� ̃�U�l$$VW�|$(;���u_^�   ]��� S�����ΈD$,�����N�^UWj �D$<�:���PjS��	 �������D$��   �N��~$9N0u�N,UWj ����PjS���	 �����D$����   ن�  ن�  ������uHل��  �\$ل��  ٜ��  �D$ٜ��  ل��  �\$ل��  ٜ��  �D$ٜ��  ن�  ن�  ������uHل��  �\$ل��  ٜ��  �D$ٜ��  ل��  �\$ل��  ٜ��  �D$ٜ��  �L$Q��D�C ��P���� ����[t<h�D����"����t,UW���������  �|$( t���X����|$, t�������D$_^]��� ������������̃�U�l$V��N2���L$��   ;���   W�ΈD$ �������|$$ttS��������ΈD$$�����؋D$;CuU���3���;l$�D$(}.�S�Lm �ʋ��W�P�O�H�W�P�O�H�W�P�W���3����|$( t�������[;l$W}�N�Dm ���������L$������T$R�N�����|$  _t���G����^]��� ������������́�   SUVW���w 3�2�;���  �L$,�����L$D�����L$����9wD}	V�O8����9oD|�o@�D$hP��D����P�����;��R  h�D���!�����>  ���������/  �������;����  �t$�w�.�C��I�ȋN�IR�ȍT$lR��������L$,�P�T$0�H�L$4�P�T$8�H�L$<�P�T$@�N�C�v�I�ȍvR�ȍT$lR��������L$D�P�T$H�H�L$L�P�T$P�H�L$T�P�D$DP�L$0�T$\Q�T$pR������L$ �P�T$$�H�L$(�P�T$,�H�L$0�P���L$�T$(�����D$P�L$`�	����L$\Q�O8�������l$�����_^]�[�Ĕ   �;��  3ۋ���I �w��G�I�N���IR����$�   R�������P�L$0������N�G�v�I���vR���T$lR������P�L$H�����D$DP�L$0Q��$�   R������L$ �P�T$$�H�L$(�P�T$,�H�L$0�P���L$�T$(�����D$P�L$`�����L$\Q�O8����������-���_^]�[�Ĕ   Ã�89ot�G;�t�UP�B���Љo�o�o_^]��[�Ĕ   �j�h�Hd�    P��(SUVW�  3�P�D$<d�    ��t$�n �~�L$02ۉl$$�|$��������  ����  �F ��~9F@u�D$����������D$�f  �L$(�+J W�L$,�D$H    ��J ��W��j V�|$,�F� ����~Z�\$$3�D$�x�L$�Q�������t/������G���O���W;W����t
�G��������u��|$ W�L$,�J �|$��3�3���~
���;�|�Q�L$,�9J ��~%�T$����+��9 t�����    ����u�3�9T$$��   �T$ �L$�AD$ �����   ;L$��   �x����   �\$;��~   �x��|w;�}s�x��|l;�}h�x;�ta�X;�tZ;�tV�x;�t	;�tK9xtF�<��\� �����H�<��\� �����H�<��\� �����H9Ht���|� �����D$ ��;T$$�:����\$�|$��(W�������{ |�C    ��~w+��|$$�L$0�W����<.��x"�M ���@�D$�H<��R�L$4�½����yލL$0�t�����u����\$�L$<���T$�$�%����D$0P���������l$$u��L$(�D$D�����I �D$�L$<d�    Y_^][��4ÊËL$<d�    Y_^][��4�U����j�h6Id�    P��h  SVW�  3�P��$x  d�    ��^3�2�;߉\$$�  9�  �s  ;�~
9^0�D$t�D$ S�N(�ї���L$L�h����L$d�_�����$�   �S�����$�   �G�����$�   �;�����$�   �/����L$|�&�����$,  ������$  �����|$,�|$0�}��Plj �L$8Q����j��Ǆ$�      诵��� �L$4�\$DǄ$�  �����e ��Plj��$�   Q����j��Ǆ$�     �n���� ��$�   �\$4Ǆ$�  �����! �F3�;���  9�l  ��  ;��q  �L$(�L$ �\$$��  D$ � �@���\$D���T$4��D��z��Dz�   ��   ���D�   {�   �D$,PS��$�   Q��$�   R��$�   P��$�   Q��$�   R�D$hP���\$���$�la �L$dQ��$�   R��$�   P��$�   Q��$�   R��$�   PS���	 ��h  �T$<���$0  Q�H��$L  RQP��$8  R��$4  P��$�   Q��$�   R��$�   P��$�   Q��$   R��$  P� 
 �\$t��L�L$LQ�N��L����|$ t�N,�T$dR��6����D$ ���l$$�\$(��������H����  8L$��   ;��  �D$$3ۉL$ �D$$��  D$ � �@���\$D���T$4��D��z��Dz�   ��   ���D�   {�   �L$,QP�T$lR�D$XP���\$���$�nn �L$LQ�N������N,�T$dR��p����D$ ���l$$�j����f;�~b�D$$�L$ 3ۉD$$���$    ��  �D�L$,Qj �T$T�R���\$��� �$�] �NL$ �D$LP�����D$ ���l$$u��F ��~9F@u�������h�   ��x  j W�蝊 ���W���W@�Whݟ�   �苆�  ��ٖ�  ٖ�  ٖ�  �hEٖ�  ٖ�  ٖ�  ٖ�  ٖ�  ٞ�  ٖ�  ٖ�  ٞ�  tP��K����ǆ�      �Ë�$x  d�    Y_^[��]� ��S�\$��UVW����   3�9~tm�^��xT��i�   ��    �F��(�    ��(�   ��Ht�G��tj P����H3��G�G�G����   ��}�3���F�RWP���҉~�~�~_^][� �F;�}y�N��PSQ����3�;FtU�N��+�iɰ   i��   WR�Q�1� �F��;�}$����i��   +�F�P���^����ǰ   ��u�_�^^][� _�V�V^][� ��   ���;�|U��+�i�   ���D$�N��)�    ��)�   ��Ht�G��tj P����H3��G�G�G��   �l$u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� �����������U������   SVW���z����ˈD$"������|$" �D$#t��t���I������D$!u�D$! �uV���`��j ���wF���\$8�|$! �{�|$4t�������D$!�'�KVj 輵��PjWj j��	 �����D$!��  ��x  W�_������u��W�D$DP���M@���    ���u�{HW��^������u��W�L$DQ���!@���    ���u���   ��~O�D$$    �D$(���   t$$V�^������u�M�~W�T$DR��?���    ���D$$�   �l$(u��u�D$8��$����D�Cz$����   9C0��   ��� �����������   ��~a9C0u\�L$@�>���D$@P����E���\$(�K,�T$@Rj 胴��P�D$<jPj���	 ���\$<�����D$!����Au��薣����������|$! �T  �C ��~9C@u���q����C���6  ��l  ;��(  �D$8��������������4����������   �������������D��   ��������D��   �F(������D��   �FP������D��   ������������������������Azu������h  t� ���Ƀ����X����H��X�u��؍��  �   ���> t$�S,��h  ����$R��l  P�RP�7�����؃���u��9�������������hT��h�Sh�  h�E�p� ���D$! ���������ٓ�  ٓ�  ٓ�  �hEٓ�  ٓ�  ٓ�  ٓ�  ٓ�  ٛ�  ٓ�  ٓ�  ٛ�  �D$8����;����Az��8  �����|$" t�������|$# t���F����D$!_^[��]� ��������j �DI�S������V��j �DI�@����D$t	V��E������^� ����������QUV�t$��;���   �FS3�;��][^��]Y� 9E}P�����9]t�F;ÉE�\$~�W����    �t$�F�U�Ӌ����&   󥋈�   ���   ���   ��   P�B�ЋD$���ð   ;E�D$|�_[^��]Y� ^��]Y� j�h&Jd�    PQSUVW�  3�P�D$d�    ��t$�@_	 3ۍN�\$ �TT�<� �F0I�^�^ �^$�N(�D$ �o� �N8�D$ �b� �~H�o���D$ �P:��h�   SW�� ���U ���W@���   �Whݟ�   �e� ǆ�   DI���   ���   ���   ��   �D$ ��� h@h`�jj��  P�D$4迩 h@h`�jj��@  Q�D$4蠩 ��`  ǆd  XI��h  ��l  ��p  ��x  �o���D$ 
�9��h�   SW�� ����U �W@�Whݟ�   ǆ  �H��  ��  ��  ǆ   �H��$  ��(  ��,  ��4  ��8  ǆ<  �$��@  ��D  ��H  ǆL  �H��P  ��T  ��X  ǆ\  �H��`  ��d  ��h  ǆl  I��p  ��t  ��x  ��|  ���  ��ݖ0  ��ݞ8  �D$ ���  ���  ���  ���  ���  ���  ���  ���  ��8  ���  ���  ���  ���  �|������  ��0  �ƋL$d�    Y_^][�������������j�hKd�    PQSUVW�  3�P�D$d�    ��t$�\	 �|$,3�W�N�\$$�TT�� �D$(;ÍN�D$ �0I�Y�Y�Y~P�����D$0�؍N(�D$ �#�P�� �N8�D$ �}� �~H�o���D$ �k7��h�   SW�� ��L$@�U ���W@���Whݟ�   �#L$,Q���   �� ǆ�   DI���   ���   ���   ��   �D$ ��� h@h`�jj��  R�D$4�ͦ h@h`�jj��@  P�D$4讦 ��`  ǆd  XI��h  ��l  ��p  ��x  �o���D$ 
�6��h�   SW�& ����U �W@�Whݟ�   ǆ  �H��  ��  ��  ǆ   �H��$  ��(  ��,  ��4  ��8  ǆ<  �$��@  ��D  ��H  ǆL  �H��P  ��T  ��X  ǆ\  �H��`  ��d  ��h  ǆl  I��p  ��t  ��x  ��|  ���  ��ݖ0  ��ݞ8  �D$ ���  ���  ���  ���  ���  ���  ���  ���  ��8  ���  ���  ���  ���  �������  ��0  �ƋL$d�    Y_^][��� ������SVW�������P0j����h�   3ۍ~HSW�} ���Wh�   �W@S�Whݟ�   ��x  W�w} ���W���W@�Whݟ�   9^�~t�G;�t�SP�B���Љ_�_�_9^$�~t�G;�t�SP�B���Љ_�_�_9^4�~(t�G;�t�SP�B���Љ_�_�_9^D�~8t�G;�t�SP�B���Љ_�_�_9��   ���   t�G;�t�SP�B���Љ_�_�_S���   ����9�  ��   t�G;�t�SP�B���Љ_�_�_9�p  ��d  t�G;�t�SP�B���Љ_�_�_��  9^t�F;�t�SP�B���Љ^�^�^_^[�������U����j�hKKd�    P��   SVW�  3�P��$�   d�    ���'����}3��D$X�D$T�D$TP�L$\Q���Y> �؄��I  �D$X��t	���7  3��T$HR�ωD$L�D$`�G' �؄���   �D$\P���1' �؄���   ��@  Q���)) �؄���   ��P  R���) �؄�t|��  P����( �؄�th��   Q����( �؄�tT��0  Rj����& �؄�t>���  Pj���& �؄�t(���  Qj���& �؄�t���  Rj���q& �؄��D$D����ti�D$DP���g& �؄�tW�D$D3�+�t(��t��uE���  t<Ɔ�  ���  ���  �'���  Ɔ�  tƆ�  ���  ���  �3Ʉ��D$C �L$L�L$d�L$h��   �L$CQ���#$ �؄�tr�|$C tk�T$dR�D$PP���n �؄�tT�|$L � @u;jh�9���؃���t���>n����W���  �pt�����3�W���  �^t�����2ۋ���c ��u2ۄ��D$D    �  �|$D��   �L$CQ���# �؄���   �|$C ��   3��T$d�D$L�D$d�D$hR�D$PP���Pm �؄�tl�|$L � @uSj@�	9�����D$`��Ǆ$�       t	��蜗���3��L$D����  �T$D����  WǄ$�   �����w�����2ۋ��$c ��u2ۃD$D���6����I��tE�D$\�L$HWPQ��蹇���؄�t-�D$X��uW���h�������u�T$HWR���\������2ۃ|$T|+����`  �D$Pt�L$PQ���$$ �؃|$P ��`  �|$X��  �|$T��  ���/  �FHP���& �؄��  �|$H �  �L$P3�Q�ωD$T�D$d�R
 �؄���   �L$P����   �D$H����;�ug��   P�Q]����  �T$P�L$`QPR���9Y
 �؄�t�D$HP��   �������� ����   ��  ��  PP�jQ�� ���oh�Th�Th~  h�E�͒ �����Ӑ =i/�C�D$P�u;��r6����   P�\����  �T$`RP�D$XP���X
 ��   ���+����2ۃ|$T|`���y� =:�|R��tW�NH�z���؃|$T|<��t8���  Q����  �؄�t$���  R���  �؄�t���  P���  �؃�   �-  �F���"  9��   �  ��  �q������  ��   �^�������   ��@  ��������   ��P  �؟������   �~\ ��   �FHP�D$d�M��������   �L$H��   Q���|[��� |�G    �L$t������L$l����3�9D$H�D$D~b����   ���T$l�D$l�D��T$t�L$|Q�T$x�D$t�D$tRݔ$�   ���\$�$�oh�����D$tP��������D$D��;D$H�D$D|��L$`�v����Ë�$�   d�    Y_^[��]� �����������j�h{Kd�    PQ�  3�P�D$d�    h�  ��4�����D$���D$    t�������L$d�    Y���3��L$d�    Y������������j�h�Kd�    P��SUVW�  3�P�D$d�    �ًl$,;���  �����U����P	 �EP�K�B� �S�R�K�EP�ҍE(P�K(�'� �M8Q�K8�� ���   R���   �I� ���   P���   �'�����   Q��   ��� ��   �R��   ��   P�ҋ�0  ��0  ��x  ��x  �&   �uH�{H�&   󥋍@  ��@  ��D  ��D  ��H  ��H  ��L  ��L  ��P  ��P  ��T  ��T  ��X  ��X  ��\  ��\  ��  ��  ��  ��  ��  ��  ��  ��  ��   ��   ��$  ��$  ��(  ��(  ��,  ��d  �@��,  ݅0  ݛ0  ��d  ݅8  ݛ8  ��`  ��`  ��d  R�Ћ�  �R��  ��  P�ҋ�4  ��4  ���  ��tP�4����ǃ�      ���   t'jh�d2������t���  �   ����3����  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  ���  �����  ���  +��D$,   �.��t�M0��� U�3�����    �<7 tEj@��0������l$���D$$    t�7�M0�D$�Θ���L$Q���n���3��D$$�����.���l$,u��ËL$d�    Y_^][��� ��j�h�Ld�    PQSVW�  3�P�D$d�    ��t$�TT�D$   �������8  3ۉ�D$�����9�,  ��   �D$��Ht�G;�tSP����H�_�_�_9�  ��  �D$
��Ht�G;�tSP����H�_�_�_9�p  ��d  �D$	�XIt�G;�tSP���dI�_�_�_h@jj��@  P�D$,讖 h@jj��  Q�D$,蔖 9�  ��   �D$�lIt�G;�tSP���xI�_�_�_���   S�D$ �DI�h���9��   ���   �D$��It�G;�tSP����I�_�_�_9^D�~8�D$��Jt�G;�tSP����J�_�_�_9^4�~(�D$��Jt�G;�tSP����J�_�_�_9^$�~�D$�0It�G;�tSP���<I�_�_�_9^�~�\$��Ht�G;�tSP����H�_�_�_���D$������J	 �L$d�    Y_^[���j�h�Ld�    PQVW�  3�P�D$d�    ��h�  ��-�����D$���D$    t���������3����D$����tW�������ƋL$d�    Y_^������������VW�|$��t5h8@���z�����t%�t$��th8@���b�����tW�������_�^�_2�^�������������V�������D$t	V�;/������^� ��j�h�Md�    PQSUVW�  3�P�D$d�    ��t$�@I	 3ۍN�\$ �TT�<� �F0I�^�^ �^$�N(�D$ �o� �N8�D$ �b� �~H�o���D$ �P$��h�   SW��l ���U ���W@���   �Whݟ�   �e� ǆ�   DI���   ���   ���   ��   �D$ ��� h@h`�jj��  P�D$4迓 h@h`�jj��@  Q�D$4蠓 ��`  ǆd  XI��h  ��l  ��p  ��x  �o���D$ 
�#��h�   SW�l ����U �W@�Whݟ�   ǆ  �H��  ��  ��  ǆ   �H��$  ��(  ��,  ��4  ��8  ǆ<  �$��@  ��D  ��H  ǆL  �H��P  ��T  ��X  ǆ\  �H��`  ��d  ��h  ǆl  I��p  ��t  ��x  ��|  ���  ��ݖ0  ��ݞ8  �D$ ���  ���  ���  ���  ���  ���  ���  ���  ��8  ���  ���  ���  ���  �|����T$(R�Ή��  ��0  ������ƋL$d�    Y_^][��� ������������V�t$��th�F���;�����t��^�3�^���������������̸�F�����������V��Fh`/P�A������u �D$����  hxYP�( ��3�^� �N@耥����u �D$����  hDYP�u( ��3�^� ���   ���q  �$�@(���   �% ��~ �D$���e  h YP�0( ��3�^� ���   �\����t �D$���6  h�XP�( ��3�^� ���    ��   �D$���	  hpXP��' ��3�^� �D$����   h�WP�' ��3�^� ���   �% ��t �D$����   h�WP�' ��3�^� ���   �����u �D$����   hPWP�V' ��3�^� ���   u*���   <tE<tA�D$��tXh WP�#' ��3�^� ���    t�D$��t3h�VP��& ��3�^� �   ^� �D$��thhVP��& ��3�^� �&E'e'e'V�񃾈   u>h�Yh�Yh|  h�Y苃 �����   ��# 3Ʌ����������   ��^Ë��   ^��������������̋D$��w�$��(�   ø   ø   �3�ÍI �(�(�(�(�������̸   ����������̋D$��t�A@��AH�X�AP�X�D$��t�AX��A`�X�Ah�X��@�Ƣ����� ��(�h$ ��������j�h�Md�    PV�  3�P�D$d�    ��D$P�L$��( j �L$�D$    ��1 �L$��" ��t
�N(�! ��L$Q�N(�H) �L$�D$�����! �L$d�    Y^��� ����V�t$��thpG���[�����t��^�3�^���������������̸pG�����������SU�l$VWU���B	 �E�C�M�K�U�S�E�C�u�{�    󥍵�   ���   �   �_^]��[� ���������������j�h&Nd�    PQVW�  3�P�D$d�    ��t$��A	 �~���D$    �4Z�:�����   ��� �`/�F�d/�N�h/�V�l/���D$�F�� ���ƋL$d�    Y_^����������������j�hXNd�    PQV�  3�P�D$d�    ��t$���   �D$    ��� ���D$�����A	 �L$d�    Y^�������́�   V��Fh`/P�i<������u%��$  ��th�ZP�\# ��3�^��   � �NQ�T$Rj ��$�   P�#�����~���`V���L$�$�y"����u%��$  ��t�h�ZP��" ��3�^��   � �   ^��   � �VW�|$j ��j����& ��t,�FP����" ��t�NQ���D ��t�Ƙ   V���E _��^� ����̃�VW�|$��D$P�L$Q���D$    �D$    �& ��t@�|$t2�_��^��� �VR��� ��t�FP��� ��t�Ƙ   V���P _��^��� ����̸   �����������U����j�h�Nd�    P��hSVW�  3�P�D$xd�    ��}���]tW��tS�} tTS�L$�����PW�L$4����P�L$L�o� ��Ǆ$�       �}������L$D�EǄ$�   ������ ��E    ���   �O������
  �M����   ݆�   �����z݆�   �݆�   �_����z	݆�   �_݆�   �_����z	݆�   �_݆�   �����Au݆�   �݆�   �[����Au	݆�   �[݆�   �[����A��uw݆�   �[�L$xd�    Y_^[��]� ��t݆�   �݆�   �_݆�   �_��t݆�   �݆�   �[݆�   �[�   �L$xd�    Y_^[��]� �E�L$xd�    Y_^[��]� ����́�   SU��$�   VWU����A	 �{W�D$P���W����    �U���   �b� _^]�   [�Ā   � ��������������̸XH����������̸�   ����������̋L$h�Z�% �   � ���������̸@I�����������j�h�Nd�    P��VW�  3�P�D$ d�    ��t$蠸 ���   ���D$(    �T[�e �D$P�@I�D$,�������N�P�V�H�N�P�V� 0�F�0�N�0�V �0�ωF$�F(   �* Ɔ�    �ƋL$ d�    Y_^�� ����������������j�hOd�    PQVW�  3�P�D$d�    ��t$�T[���   ���D$   � 2��ψ��   �D$� ���D$�����ڸ �L$d�    Y_^�����������VW�|$��;�t8S���   ���f W��Ɔ�    �G� ���   P����! ���   ���   [_��^� ����́��   �E ������ ����������́��   �u �   ����������������V��L$���   PjQ�zw	 ��P���   �k ^� �������VW�|$j j��h � @���� ��u_3�^� S���   P��2��, ��t���   Q���E ��t����LF ��u2���[_^� ������������̃�UV��W���   ���; �l$3��D$�D$�D$P�L$Q�Ƽ   h � @��� �nT ��u_^3�]��� S2ۃ|$uW���� ��tV���1 ��t����DH ��u2���[_^]��� ́��   �� ������������������̋L$h�[�! �   � ����������S�\$��U��~[W�|$��|QV�t$��|G;�tC�E�;�9;�5�M�;�~�;�}��P����B���E����S����WV��] ��^_][� ����VW�|$��;~tdS3�;�~C9~~�~�N��PWQ����;ÉFt9�N;�~��+���R��SP�] ��[�~_^� �F;�t�SP�B�Љ^�^�^[_^� ����������S�\$��V��~[U�l$��|QW�|$��|G;�tC�F�+;�9;�5�N�;�~�;�}��P���6����F��    R��Q��R��\ ��_]^[� ����SU�l$VWU���8	 �C�@�K�UR�ЋM�K�U�S�E �C �M$�U(�K$R�K(�} �E,P�K,�q �M0Q�K0�e �U4R�K4�Y �E8�C8�u@�{@�   �Mp�Kp���   �ExR���   �[x�( ���   ���   ���   ���   ���   R���   �� ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   �   �_^]��[� VW�|$��t5h�F���������t%�t$��th�F���������tW������_�^�_2�^�������������VW���������G�����   �O(�� �O,�� �O0��� �O4��� ���   ��� _�^����������������j�h;Od�    PQ�  3�P�D$d�    h�   �5�����D$���D$    t���;����L$d�    Y���3��L$d�    Y������������j�hkOd�    PQVW�  3�P�D$d�    ��h�   �������D$���D$    t����������3����D$����tW���M����ƋL$d�    Y_^������������VW�|$��t5hpG���J�����t%�t$��thpG���2�����tW�������_�^�_2�^�������������V��������D$t	V�������^� �̋D$VW��3�9��   ~&���   ���   �Q�RP�vq	 ����;��   |�_^� ���VW�|$jj��h � @���� ��u_3�^� ���   ���   SPQ��2���� ��t6���    ���D$�D$P�? ��t8\$t���   Q����� ��t����$@ ��u2���[_^� �����3�9��   �������j�h�Od�    PQ�  3�P�D$d�    h�   �������D$���D$    t�������L$d�    Y���3��L$d�    Y������������j�h�Od�    PQVW�  3�P�D$d�    ��h�   ������D$���D$    t���������3����D$����tW��������ƋL$d�    Y_^������������VW�|$��t5h@I���
�����t%�t$��th@I���������tW���v���_�^�_2�^�������������j�h�Od�    P��VW�  3�P�D$ d�    �D$P�@I������|$0P����������th@I���~�����uB3�8D$4t<h�   �x�����D$���D$(    t���������3�V���D$,���������ƋL$ d�    Y_^�� �����V���(����D$t	V�������^� ��V��~ ��[t%�F��tj P��[�F    �F    �F    ^�����������V��L$��|3�F;�},+���P�APQ���,����F��F3���F��H�H�H^� ��������������j�h(Pd�    PQVW�  3�P�D$d�    ���L$�2 �t$ ���D$    t.V�L$�H j �L$�M  �L$�t ����t
f�> u3�����PW�*���������t'��u��Bj�����V���   �� �L$$���   �L$�D$������ �L$d�    Y_^��� ����̃�VW�D$��P�@I�����P���r�������t?h@I���p�����t/���   �� ��t f�8 t�|$P���k ���   �T$ �
��|$���B �D$ �  ���T ��_^������ �����V��~ ��[t%�F��tj P��[�F    �F    �F    �D$t	V��������^� ������V��~ �\t%�F��tj P�\�F    �F    �F    ^�����������V��L$��|*�F;�}#+���P�APQ��������F��F�N��    ^� �������V��~ �\t%�F��tj P�\�F    �F    �F    �D$t	V�������^� ������j�h�Pd�    PQSVW�  3�P�D$d�    ��t$�/	 3��\�\$�F�[�^�^�^�N(�D$� �N,�D$�{ �N0�D$�n �N4�D$�a �N@�D$�� �~p���D$��R ���   �D$�5 ���   �D$������`/�F�d/�N�h/�V �l/�^x���   �D$	�F$���   ���   ��  ���   �^8���   ���   ���   �ƋL$d�    Y_^[���j�hCQd�    PQSVW�  3�P�D$d�    ��t$�\���   �D$   �M������   �D$�} �Np�D$�PR �N@�D$�C� �N4�D$�V �N0�D$�I �N,�D$�< �N(�D$�/ 3�9^�~�\$��[t�G;�tSP����[�_�_�_���D$�����-	 �L$d�    Y_^[������������������j�hhQd�    PQSUVW�  3�P�D$d�    ���O(�� 3�;�u��7�t$(Phx^V�6 hp^V�+ ���   ����w9�$��Bhd^�0���   �D ��~h^�h�]�h�]�h\]�hP]V�� ��h�&V�� hH]V�� ���GP��� h�&V� ���O,�< ;�tf9tPh4]V� ���O0� ;�tf9tPh(]V�g ���O4�� ;�tf9tPh]V�G ��V�Op�Q ���   �� h]V���# ��;���   f9] ��   ���   :ø�\u��\PUh�\V�� �����c �L$�
 �L$(Q�T$R�ω\$(�\$0�a�����t7�L$�T ;�tf9u��78\$(��\u��\QPh�\V� �����   Ph�\V�t h�\V�i ��V���   �:������ �L$�D$ �����	 �h�\V�5 ���oUh�\V�# ��;�~l��� �OQ���j h�&V�� ����~hdRV�� ���0��~+�   ����W�R���- h�&V�� ������u݋��p V�O@�w����L$d�    Y_^][��� ��?@@%@j�h�Qd�    P��SUVW�  3�P�D$(d�    ���t$8jj���H �؄���   �GP���c �؄���   ���� ��|D���   u;3��D$�[�D$�D$ �D$$�L$Q�ΉD$4�2 �L$���D$0����������WR����1 �؄�tQ�G(P��� �؄�t@�O,Q��� �؄�t/�W0R��� �؄�t�G4P���z �؄�t�O@Q����- �؋������ۋ�l$�  U���	 �؄���   ��u2�L$8�s �T$8R���D$4   � �L$8���D$0�����l ����   P���� �؄���   ��Vu��9��������   �v����؄���   �Op�opQ���	 �؄�ts�Gx�����$�
 �؄�t]�|$ u�D$ �
���   �T$�D$P���3 �؄�t3V���M �؄�t%���   Q��� �؄�t���   R��� ���ËL$(d�    Y_^][�� � ������������V�񍎐   �r ���   �'���3�PP�Έ��   ���   ���   ���   �����^���SVW��3�3�9��   ~*���   ��;�t	��Bj�Ћ��   ����;��   |�9��   ���   t�G;�t�SP�B���Љ_�_�_���   ;�t��Bj�Љ��   _���   ^[�Ŵ �����j�h�Qd�    P��UVW�  3�P�D$$d�    ��t$�� 3퍾�   ��^�l$,�\�o�o�o���   �D$,�n� �D$P�XH�D$0������N�P�V�H�N�P�V� 0�F�0�N�0�V �0�F$�F(   9ot�G;�t�UP�B���Љo�o�o���   �ƋL$$d�    Y_^]�� ����������������j�h$Rd�    PQSVW�  3�P�D$d�    ���|$��^�D$   �3������   �D$�� 3�9��   ���   �\$�\t�F;�tSP���\�^�^�^���D$�����`� �L$d�    Y_^[���������������̃�SVW�������|$ �D$P�L$Q3�h � @�ω\$ �\$$�/? ��u_^3�[��� �|$�\$ ��   ���   R���� ��tr9\$~g�D$P�ψ\$�� ��tX8\$tM�L$Q�ω\$�� ���L$u;�t��Bj���+Q�#����;É��   u�L$;�t��Bj����D$ ���2 ��t�\$ _^��[��� ��j�hKRd�    PQ�  3�P�D$d�    h�   �������D$���D$    t��������L$d�    Y���3��L$d�    Y������������j�h{Rd�    PQVW�  3�P�D$d�    ��h�   �q�����D$���D$    t���W������3����D$����tW�������ƋL$d�    Y_^������������V���H����D$t	V�	������^� �̃���UV��W�^x3��nx���   �|$�|$Ɔ�    �� ���   �~pƆ�    � �|$ �D$P�L$Q���z	 ���@  �|$St2��s�VR���� �؄�tb�FP���� �؄�tQ�N(Q���I� �؄�t@�V,R���8� �؄�t/�F0P���'� �؄�t�N4Q���� �؄�t�V@R���� �؄ۋ��   �D$$t5�L$$Q����� �؄�t#�T$$R�I������   �����   P����� �؃|$|��tW���   �����؃|$��   ���D$    t�D$P���� �؋L$Q�� �����Fpt��tjP��� �����|$�] ��   ����   U����� �؄�t{���   P���� �؄�tg�|$|`W�Np�"F �؄�tQ�|$|J���   R���� �؄�t6�|$|/�D$P���D$     ��� �؋D$��t�H����   w���   ���   u"���   �  ��~ǆ�      ����0������   u1���   <r<v����� ��2�����   ��[_^]��� ��[_Ɔ�    ^]��� _^��]��� ������j�h�Rd�    PQ�  3�P�D$d�    h�   �%�����D$���D$    t���[����L$d�    Y���3��L$d�    Y������������V���(����D$t	V��������^� ��j�h�Rd�    PQVW�  3�P�D$d�    ��t$�|$ W�-����\8�O�N�W�V�O�N�W�V�O�N�W�V�O �N �W$�V$�O(�N(�W,�V,�O0�N03��N4�W4R�D$�H8�A�A�A�T:���GD�FD�OH�NH�WL�VL�GP�FP�OT�NT�WX�VX�G\�Oh�F\�G`Q�^`�Nh�D$�
 �Wl�Vl�Gm�Fm�On�Nn�Wo�Vo�ƋL$d�    Y_^��� ���j�hSd�    PQSUVW�  3�P�D$d�    ���|$�\$(���   9��   ���   }P���U������   3���~c���$    ���   �<���t>jp�<�����D$(���D$     t
W���a����3��L$(Q���D$$�����D$,�% ��;��   |��|$���    t:jp�������D$(���D$    t���   R�������3��D$ �������   ���   ���   S���� ����� �L$d�    Y_^][��� ��j�hKSd�    PQVW�  3�P�D$d�    ��h�   �Q�����D$���D$    t���������3����D$����t;�t�������W���� W���Z����ƋL$d�    Y_^���������VW�|$��tHhXH���������t8�t$��t0hXH��������t ;�t���s���W��蛙 W�������_�^�_2�^����������j�h�Sd�    P��TSUVW�  3�P�D$hd�    �\$|�l$xSj���'D ��t$�����������t$}(��thaS��� ��2��L$hd�    Y_^][��`ËE �P4���҃���   �E �P4���҃�t3��t�E �P4����Ph�`S�� ��2��L$hd�    Y_^][��`ÍD$8P���� 	 �L$8�D$p    �G{����u9��th�`S�D� ���L$8�D$p�����`� 2��L$hd�    Y_^][��`��D$H����������DzA�D$`������Dz6�L$8�D$p������ ��t~3���U��L$hd�    Y_^][��`��؅�th�`S�� ���L$8�D$p�����ӵ 2��L$hd�    Y_^][��`Ë\$|W����0 ����t}����   ���Ѕ���   W�L$,Q����0 �؋�Rh�D$P���D$t   ��S���D$t��|���L$���D$p�U� �L$(�D$p�����D� ��ul��;|$�v���� ������l���Wh``S��� ��2��L$hd�    Y_^][��`Å��?���Wh4`S�� ��2��L$hd�    Y_^][��`ËD$|��tWWh�_P�� ��2��L$hd�    Y_^][��`�������U����j�h�Sd�    P��(  SVW�  3�P��$8  d�    �uX��t��������]\��t��������M �u����u$�M ��s����u2���$8  d�    Y_^[��]ÍM8�zu����u�M8��s����t�����T$�L$t�T$�$�m���EP��t7� �L$\�\$\�@�\$d�@�\$l�-u����u�L$\�s����u	�L$\�n����$�   ��= �E�M�U��$�   �E��$�   �M��$�   �U��$�   �E ��$�   �M$��$�   �U(��$�   �E,��$�   �M0��$�   �U4��$�   �E8��$�   �M<��$�   �U@��$�   �ED��$�   �MH��$�   �UL��$�   �E ��$�   P�M8��$�   Q�T$LRǄ$L      ��t�����$�   �P��$�   �H��$�   �P��$�   �H��$�   �P����$�   ��$�   ��s����u��$�   �<r����$�   ��= �}T��$�   PhhY���i����t���    ���}T�uX��_�\$l�����   �L$\�s������  �D$l��ݜ$�   �L$\���\$�D$t�\$�D$|���$�k���L$D�t������  �L$D�Vq���T$|���$�b��������  �L$D�sq�����|  �����$  �$��������D$t�����D$L��������ݜ$  �D$D����������ݔ$  ݜ$$  ����ݜ$,  ݔ$T  ݜ$|  t�}X�    ��$  �}T��$�  ������D$t��=��=���ĉ� >�P�>�H�>�P�>�H�L$\�P�T$`���ĉ�L$|�P��$�   �H��$�   �P��$�   �H���P�\$݄$�   ��$�  �$�o�����t%��$�  P��$  Q�������    �����}T��$  R��$  P��$�  Q��$�  R���_������X����    ��󥍌$�   Ǆ$@  ������ ���$8  d�    Y_^[��]�S�N��j���N ��j�����^8�NH���^@��j��3ۍNp�^`�^d�^h�^i�^j�^k�j�����   �j����ݞ�   ���   ��[ݞ�   ���������������U�l$;��Q  �Kd��t��Pj���Cd    VW�u�{�   �E8�C8�M<�K<�U@�S@�ED�CD�MH�KH�UL�SL�EP�CP�MT�KT�UX�SX�E\�C\�M`�K`�}d _^t�Md��Bd���3��Cd�Mh�Kh�Ui�Si�Ej�Cj�Mk�Kk�Up�Sp�Et�Ct�Mx�Kx�U|�S|���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ]�SV��3�8^jWt?�~p���zo����t1��_ܞ�   ����z�������Dz�^x����D{	��ػ   �~k tJ���   ���2o����t9��_ܞ�   ����z&�������Dzܞ�   ����D{_��^��[��؃�_^��[����������������V��~h u�~i t"�F`��|�Nd��t��u����   �҅�u03�^�~*Q��
 ����t�j ���S( ��t���ȋ��   �Ѕ�tЀ~h t3�8Fi^���D ø   ^�����U������4  SV��W�D$�~P����	 �E��$����D��   �~j ��t�^p�3��F8���L$0�$Q���x�	 �Uj �NH�1j RS���ԉ2�q�r�q�r�q�r�q�I�r�J�T$8���̉�T$T�Q�T$X�Q�T$\�Q�T$`�Q�T$d�Q����̉�P�Q�P�Q�P�Q�P�@�Q�A�{�����X_^[��]� ��$����Dz�~k t�F@���   �4����F@3��*����L$@������$�   �����~j t�^p�3��F8���L$0�$Q���}�	 j j �T$HR�VHS���̉�VL�Q�VP�Q�VT�Q�VX�Q�V\�Q�T$8���̉�T$T�Q�T$X�Q�T$\�Q�T$`�Q�T$d�Q����̉�P�Q�P�Q�P�Q�P�@�Q�A������X��u2�_^[��]� �~k t���   �3��F@���L$0�$Q����	 j j ��$�   R�VHS���̉�VL�Q�VP�Q�VT�Q�VX�Q�V\�Q�T$8���̉�T$T�Q�T$X�Q�T$\�Q�T$`�Q�T$d�Q����̉�P�Q�P�Q�P�Q�P�@�Q�A������X���6�����E�E���D$@��݄$�   ������D$H��݄$�   �����X�D$P��݄$�   �����X�D$X��݄$�   �����X�D$`��݄$�   �����X �D$h��݄$�   �����X(�D$p��݄$�   �����X0�D$x��݄$�   �����X8݄$�   ��݄$   �����X@݄$�   ��݄$  �����XH݄$�   ��݄$  �����XP݄$�   ��݄$  �����XX݄$�   ��݄$   �����X`_݄$�   ^��[݄$  �����Xh݄$�   ��݄$$  �����Xp݄$�   ��܌$,  ���Xx���]� ������W���`3�_ËGdVP�Y ������t���y}��9G`u��^_�^3�_�����������W���Gd��u_�V�w`��|~ P� ����t�w`���2}��;�t^3�_Ë�^_����̸0J�����������j�hTd�    PQSUVW�  3�P�D$d�    �ى\$�l$(U�� 3��K�t$ �4a��	 �K8�D$ �Y���KH�D$ �M`���sd�sp�   �����9`������y񍋠   ��X��U�D$$�+������ËL$d�    Y_^][��� j�h\Td�    PQV�  3�P�D$d�    ��t$�4a�Nd���D$   t	��Pj�ҍ��   �D$�J� �N8�D$�=� �N�D$ �0� ���D$������� �L$d�    Y^���VW�|$��;�tC�Nd��t��Pj���Fd    S�������P0j���ҋ�蕺��W��� W���5�����[_��^� ���������̅�t��t�8 tPhbQ�g� ������V��~d W�|$t�Nd��P0W��W���O� _^� ����������U������4SV��N`��W}/�E���Y  h8ehbP��� ����H ��_^[��]� �Fd��u/�E���#  h$ehbP��� ����H ��_^[��]� ����   P�f �؃���u/�E����  h�dhbP�� ���zH ��_^[��]� ���Wz��9F`t�M��d�  �}WS��������u
�td�}  3�9~`~'�I W���x  ��tY��ȋ��   �Ѕ�tV��;~`|܋}�^���o�	 ����   ���9  h\dhbW��� ����G ��_^[��]� �M�d�  �M��c��  �}�ȋ�BW�Ѕ�u�����  h�chbW�� ���G ��_^[��]� S�L$,Q�N ��^���L$(�d���T$ ���$�nU��������  ���D$ ��������A�j  ���$�CU�������1  ��;�\$ �����  �L$(��c�����  �L$(�ye������   �F8��$������   �F@�^8����A��   ���^@������   �^H���2e����u
��c��   �T$(R���H^������4����Au
�hc�   �~j t0�Np��d����u
�Hc�   ��_ܞ�   ����{�c�|�~k t0���   �d����u��b�`��_ܞ�   ����{��b�F�   _^[��]� �|b�1�`b�*��t-h$bW��� ����E ��_^[��]� �ظb���6����E _^��[��]� ����̃yd ��   t�Id��P���   ������V��~d t�Nd��T$�@R����D$�NQj0P�FD	 �V8RjP�:D	 �NHQjP�.D	 �VjRjP�"D	 �NkQjP�D	 �VpRjP�
D	 ��H���   QjP��C	 ���   RjP��C	 ���   QjP��C	 �V`RjP��C	 �NhQjP��C	 �ViRjP�C	 ��H�~d t�Nd�^�D$�B��^� ����������V�t$Wjj��h � @���H� ��u_3�^� �GdSP���1� �؄���   �OQ���� �؄���   �W8R���� �؄���   �GHP���R� �؄���   �OjQ��� �؄���   �WkR��� �؄�t�GpP���� �؄�tn���   Q���� �؄�tZ���   R���M �؄�tF���   P���8 �؄�t1�O`Q����� �؄�t �WhR��� �؄�t�GiP��� �؋�� ��u2���[_^� ����������̃�UV��Nd3�;�Wt��Pj�҉nd�n�����P0j���ҋ������|$�D$P�L$Qh � @�ωl$�l$� ��u_^3�]��� �|$S�Ä���  �T$R�ωl$ �:� ���Ä���  �D$;�t(P������;ŉFdu�L$;�t	��Pj��2��Z  �FP����� �؄��E  �N8Q����� �؄��0  �VHR���� �؄��  �FjP����� �؄��  �NkQ����� �؄���   �VpR���H� �؄���   ���   P���0� �؄���   ���   Q���H� �؄���   ���   R���� �؄���   3�9Fd�n`���|$�E |7U����� �؄�tq�|$|)�NhQ���A� �؄�tY�ViR���0� �؄�tH�|$}A�m ��u�Fd���|0��������t%j ��� ��t��ȋ��   �Ѕ�t�Fi�Fh���� ��u2���[_^]��� �������̸   @�����������U������x  VW�t$(�   ���V������y����S�;�[(��C�K�S�s�|$(�{�|$,�D$@�C�L$D�\$@�K����|$0���|$4���|$8���|$<�{�|$p�{�|$t�\$p�{ �|$x�{$�|$|�{(��$�   �{,��$�   �{�|$X�{�|$\�{ �|$`�{$�|$d�{(�|$h�{,�|$l�;��$�   �{��$�   ����$�   ����$�   ����$�   ����$�   �|$@�D$H�L$L�T$P��$�   �|$D��$�   �C��$�   �K ��$�   �S�t$T��$�   ��$�   ��$�   ��$�   ��$�   �K,�S$�C(��$�   �L$x��$�   �T$p��$�   �D$t��$�   ��$�   ��$�   �T$|��$�   ��$�   ��$�   ��$�  ��$�   ��$�   �$�����u��$�  R�����$�J�����u2�_^��]Í�$   ������荄$   P�����$������tыu��tb������$�1�����uO��$�  Q��$  R��������    ��$�  󥍄$   P��$  Q�M������    ����$   �T$(R��$�   P��$�  ������L$(�P�T$,�H�L$0�P�T$4�H�L$8�P�D$@P��$�   Q��$�  �T$D�c�����T$@�H�L$D�P�T$H�H�L$L�P�T$P�@�L$XQ��$�   R��$�  �D$\�!�����L$X�P�T$\�H�L$`�P�T$d�H�L$h�P�D$pP��$�   Q��$�  �T$t�������T$p�H�L$t�P�T$x�H�L$|�P��$�   �@��$�   Q��$�   R��$  ��$�   �������$�   �P��$�   �H��$�   �P��$�   �H��$�   �P��$�   P��$�   Q��$  ��$�   �=������$�   �H��$�   �P��$�   �H��$�   �P��$�   �@��$�   Q��$�   R��$  ��$�   ��������$�   �P��$�   �H��$�   �P��$�   �H��$�   �P��$�   P��$�   Q��$  ��$�   �������$�   �H��$�   �P��$�   �H��$�   �Pj �L$,Qjj��$�   �@j j�ˉ�$�   �n� _�^��]�������U����j�h�Td�    P��hSVW�  3�P�D$xd�    ��3ۍN�\$�$�	 ����  9^d��  �L$�*� �Nd��@<SS�T$R��$�   �Є��F  SV�\$�_��������0  �} �u�}�D$��   ��������   �F�_������   �F�_������   ����$�1I��������   �F���$�I��������   �F���$��H������tx�D$�����z�����D$�W����z�_����D$$�W����z�_����D$,�����Au�����D$4�V����Au�^����D$<�V����Au/�^�,�D$��D$�_�D$$�_�D$,��D$4�^�D$<�^��؍L$Ǆ$�   �����P� �D$�L$xd�    Y_^[��]� �ËL$xd�    Y_^[��]� ��������������j�h�Td�    P��4SVW�  3�P�D$Dd�    ��3ۍN�\$��	 ��t{9^dtv�L$�(� �Nd��@<SS�T$R�\$X�Є�tC�L$\QV�\$�`�������t)�|$X t�L$T��R�֙ ��|$T�   �t$��D$�\$�L$�D$L�����[� �ËL$Dd�    Y_^[��@� ����U�������4SVW�}�����$���P�����t	�_^[��]�����G(��������Dz�G ��$����Dz2����~`��   �FdP�h� ��������   ���j��9F`��   ���D$/t	��BL���Ћ�3��`j�����[  S��� ����tY��E�RDP���҅�u�D$/�B�} t<�D$0P�L$<Q��������t'����   �����D$0��Bl���\$���D$H�$�Ћσ���i��;�|��D$/_^[��]Ë}��ty�Nd��BH�Є�uk��Ndj ���$j ���������tA�NdQ��������E�RDP���҅�t�Nd���D$/t	��Pj�҉~d�/��Pj�����D$/ �D$/_^[��]ËNd��PDW�҅�t��D$/�} tA�D$8P�L$4Q�Nd������t+�Nd����   ���D$8�vd��Bl���\$���D$@�$�ЊD$/_^[��]���U����j�h�Td�    P��  SVW�  3�P��$�  d�    ���|$`�w�Ή�$,  �'�	 ����  �_H�ˉ\$X�1U������  �`�v  ��$�  P���`�	 ��$�  Q��$�   SR�U������$�   ��T����u��$�   �;S�����*  �]j���g���� ��$����Dz7j���O����@��$����Dzj���6����@��$�D$?����D{�D$? h��jj��$  P�֛��h��jj��$   Q�������F�N��$�  �V��$   �F��$  �N��$  �W ��$  �G$��$  �O(��$  �W,��$  �G0��$  �O4��$   ��$�  ��$$  R��$�   ��$,  P���r������$�   �P��$�   �H��$�   �P��$   �H��$  �P��$  P��$�   Q�ˉ�$  � ������$  �H��$  �P��$  �H��$  �P��$  �@��$�   ��$   ��S�����x  ��$  ��S�����d  �|$? t.��$�  Q��$�   R��$  ��K��P��$�  P���:������$�   Q��$�  R��$  �K�����$l  �P��$p  �H��$t  �P��$x  �H��$|  �P��$l  ��$�  ��P������  ��$  P��$  ��`���\$L��$�  Q��$�   ��`���\$L�D$D   ����At�D$D    �t$D�4v�����4�  ��4  ��4   ��$�  ��4  ��$�  ��4  ��$�  ��4�   ��$�  ��4  ��$�  ��4�   ��$�  ��4   ��$�  ��4�   ��$�  ��4  ��$�  ��$�  ��4  ��$�  ��$�  R��$p  ��$�  �J�������%�$����4����Az*���D$>������A�&  ��$�   P��$�  �M������D$> ��$l  ��L$|�P��$�   �H��$�   �P��$�   �H��$�   �P��$  P��$�   ��$�   �P_���T$L�|$> �  �|$D t���L$|Q����$�   �$R�0J����P��$@  P��$�  �HI����$  ��$<  +�R�L$H��^���D$L��4������uM�D$D��$<  ��$@  ���$D  �P��$H  �H��$L  �P��$P  �H�P�f��$�  �������$l  ��$p  ��$t  �D$|��$x  ��$�   ��$|  ��$�   ��$�  �D$> ��$�   ��$�   ��$�   ��؍�$�   P��$�   Q��$�  �XH��P��$�  R���(����t$XV��$�   P��$�  �/H��P��$�  Q��������|$? tV��$�   R���������$�  P��$�  Q��$�  �H�����$|  �P��$�  �p��$�  �X��$�  �X��$�  �@��$�   ��$�  ��$�   ��$�   ��$�  ��$�   ��$�   ��$�   ��$�   �M������  �D$|��PQ��$�  �G������$�   �$R�H����P��$8  P��$�  �[G����$4  �L������  �t$XV��$8  �fG�������%�$����4����Az"��������A��  ��$�   Q����I�����2ۍ�$4  �ۋ�T$d�H�L$h�P�T$l�H�L$p�P�T$t�@�D$xt}�|$> uv�L$|Q�L$h��F����T$|�\$LR��$8  ��F�����\$L����zD��$4  ��$8  ��$<  �D$d��$@  �L$h��$D  �T$l��$H  2ۉD$p�L$t�T$x�D$|P�L$hQ��$�   R�M������$�   �K�����o  ��$�   P��$�   �4F���|$> t��u�����%�$����4����A��   ��������AuX��$�   Q��$�   �H�����$�   �H��$�   �P��$�   �H��$�   �P��$�   �@��$�   �_��������$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��؍�$�   Q�L$h�@E��������������4��������AuJ�T$d�ڋD$h�؋L$l�؉�$�   �T$p��$�   �D$t��$�   �L$x��$�   ��$�   ��$�   �[������������zL��$�   R�L$h�G�����$�   �P��$�   �H��$�   �P��$�   �H��$�   �P��$�   �|$? t��$�   P��$�   Q�M�������$�  R��$�  P��$�  �D�����$�  �P��$�  �H��$�  �P��$�  �H��$�  �P��$�   ��PQ��$�  ��$�  ��C������$�   �$R�ND����P��$(  P��$�  �C����$$  ��H������
  ��$$  Q��$�   �C��������������4��������Au\��$�   �ڋ�$�   �؋�$�   �؉�$$  ��$�   ��$(  ��$�   ��$,  ��$�   ��$0  ��$4  ��$8  �^������������zO��$�   R��$�   ��E�����$$  �P��$(  �H��$,  �P��$0  �H��$4  �P��$8  ��$�   P��$(  Q��$�  R�J������$�  �mI����u��$�  �G������	  �D$|P��$�  �tB����$����z��$$  �kG����$�  �_G����$�  Q��$�   �;B������$�  �$R�L$p�$B�����\$��$�  ���$�@����_݄$�  ��������A��4u������Au݄$�  ����������  ����������\$��$�  �D$V �T$�$�8J���L$|��$�   ��$�   ��$�  ��$�   ��$�  ��$�   ��$�  ��$�   ��$�  ��$�  ��$�  ��=��=�5�=��=��=��$\  ��=��$P  ��$`  ��$h  ��=��$x  3ۉ�$X  ��$p  ��$L  ��$T  ��$d  ��$l  ��$t  �D$@ �D$A �D$\ �D$] �\$D�wp�T$D�D$`�|j �J  ��V�F��L  ��N�W�V�G�F�O�W�G�D$D��$T  �D@�D\�7>���|$> �W  ����\$��$T  ����\$�F�$��>����$<  �]E����$<  Q��$�  VR�wG��݄$X  ����$�  P����$�  �$Q�b@��݄$T  ��P�D$\��$�  RP����$�  �$Q�7@��݄$T  ��P��$�  R��$�   P����$x  �$Q�	@�������/?�����(?��� ݜ$<  ��$�  �@Rݜ$H  ���@��$h  ݜ$X  ݄$�  �$P�?��݄$�  �T$h��P��$x  QR����$�  �$P�?��݄$�  ��P��$�  Q��$�   R����$�  �$P�`?�������>�����>��� ݜ$�  ��$<  �@Q�Mݜ$�  �@��$�   Rݜ$�  �������$�  P��$�  Q�M�������$�   �vC���\$L��$�  �fC���D$L�����������Xe������z��$�   �}C����$�  �qC����$�  R��$�   P��$d  Q�E�����$`  �H��$d  �P��$h  �H��$l  �P��$p  �@����$h  �   �������������T$L��4������za��������uX��$�  ��P��$�   �=���\$D���d$L�B	 ݔ$�  ���\$D����Au��ݜ$�  ݄$�  ���݄$�  �������4����Az	��ݜ$�  ��$�  �D�����h�����ܔ$�  ����Dzܔ$�  ����D�H������D$>�����F��$�  Q����$h  �$R�W=���F�L$h��P��$�   PQ����$�  �$R�0=�����P��$�  P��$�   Q����$�  �$R�=�������-<�����&<����$�   P��$`  Q��  �
<���MP��$�  R������|$? t��$�   P��$`  Q�M�j�������   R��$x  P��$�  ��;�����$T  �P��$X  �H��$\  �P��$`  �H��$d  �P��$h  ��$T  �A�����m  ��$T  P��$�   �;�����$T  Q�L$h�;��ݜT  ��$T  R��$�   �;��ݔ\  ��������Au���@�����@�����L$Du�D@�����4��������u���݄T  ��������Az	��ݜT  ��_ܜ\  ����At:��4ܜ\  ����A{&���������Az"݄T  ��������Az�D@ ����D@ ��؀|@ u,��=��=��=���=�O��=�W��=�6V���:���%�$����'����Az"��N�V��F�O�N�W�V�G�O�W�D$D������0����������$�  �$������$|  �?���\$D�|$> ��  ��$�  P��$(  �	:���\$L�D$D���$�V0�������  �D$D��$����D��   �D$L���$�'0��������   �D$L������������D��   �D$D������������4����Az�������ݔ$  �������Pe���������0'u�����������������Az�������ݔ$�  �������������T$D������������Az-������������z������ݔ$�  �@������ݔ$�  �1��������������Az����3���$�  d�    Y_^[��]� ���Ƀ��T$T�$�/������t��D$L��$����D{���$�  Q��$�   �8�������\$D����Az����ݜ$�  ��  ��$�  � ��$�  ��$�  ��$�  ��$�  ��$�  ��$�  ��$�  ��$�  ��$�  ��$  ��$�   ��$   ��$�   ��$  ��$�   ��$  ��$�   ��$  ��$�   ��$  ��$�   ��$  �D$X��$  ���$   �H��$$  �P��$(  �H��$,  �P�@��$0  ��$�  ��$4  ��$�  ��$8  ��$�  ��$<  ��$�  ��$@  ��$�  ��$D  ��$�  ��$H  ��$�  Ǆ$�      ��$L  ��$P  �� ��$t  � ��$�  ��$�  ��$�  ��$t  ��$�  ��$x  ��$�  ��$|  ��$�  ��$�  ��$�   ��$�  ��$�   ��$�  ��$�   ��$�  ��$�   ��$�  ��$�   Ƅ$�  ��$�  ��$�  ��$�  ��$�   �L$d�T$h��$�  �D$l��$�  �L$p��$�  �T$t��$�  �D$x��$�  �L$|��$�  ��$�   ��$�  ��$�   ��$�  ��$�   ��$�  ��$�   ��$�  ��$�   ��$�  ��$t  ��$�  ��$�  � ��$  �̻����$�  �������$  贻����$�  註����$�  Qh�Z��$  �������$t  R��$�  ����h�Z��$x  P��$  �����E��$  Q��$�  RP��$  Q��$�  R��$  P��$  芼����胼�����|�����    ����$�  �ݔ$�  ݔ$  ݔ$  ݔ$$  ��ݔ$,  ݔ$T  ��ݔ$4  ݔ$<  ݔ$D  ݔ$L  �Pe�D$D������Aus������������Aud��4��݄$�  ����������zF��ݔ$�  ݄$  ������������z����ݜ$  �������������z��ݜ$  ������0'3�3Ƀ�tE�݄��  ����  ������������Az
��������������������A�O  ������˃���|�����|��ٍ�$t  ��Ƅ$�   ������x ��$�  Ǆ$�  ������x �M�t$`Q��蒍����$,  ��$�   ��$�   ���$�   �H��$   �P��$  �H��$  �P��$  �H��$  ��$  �V ��$  �F$��$  �N(��$   �V,�T$d�F0�D$X��T$l�N4�L$h�H�L$p�P�T$t�H�L$x�P�H�D$`3���$L  ��p��$    �|<\ tD��K��S�N�K�V�S�N�K�V�T<@�N�Tj�c����������A�����������|$> t$݄$�  �݄$�  �^݄$�  �^�Dj� ����T$���T$�$�:���D$`�Dj ���������X��������$�  �$脾����t�   ��$�  d�    Y_^[��]� j��$�  �%����@j �\$P��$�  ����� �L$Lj ��$�  ݜ$0  ������@j��$�  �\$P����� �L$L�D$Dܬ$,  ��$����{�D$D �L$D�D$`Q��$�  R�f���������$�  d�    Y_^[��]� ��������j�h;Ud�    P��   VW�  3�P��$�   d�    ��D$lP�� �L$<Q��$�   Ǆ$�       �m� �L$Ƅ$�   �|u �T$<R�D$pP�L$Ƅ$�   �Az ���   �   �t$�L$Ƅ$�   ��u �L$<Ƅ$�    ��u �L$lǄ$�   �����u ��$�   d�    Y_^�Ĝ   � V��NW3�;�t�~��Pj�҉~�N;�t��Pj�҉~�NX;�t��Pj�҉~X�N\;�t��Pj�҉~\j`WV��
 ��_^�������������SVj`3ۋ�SV��
 ����   ����^�^�^�^<�^8�^\�^X�F�F�F$�F �F�F�F4�F0�F,�F(�ND�N@�FL�FH�FT�FP^[��������������D$SV���$��2��%��������   �D$���$�%������tw�D$�D$������zb�L$3�8��   ��;�u!�����\$���   �$�_7���^��[� �   +�;�u#�Nd�ɋ�Pl���\$�$�҅���^��[� ����^��[� �����������j�h�Ud�    P��$SV�  3�P�D$0d�    �T$D3�3��\$8��   ��;�u���   �6�   ��+�;�u�yd t�Id��@h�T$ R�Љ\$8��L$�$���   ��t$@��P�V�H�N�P�V����t����L$�\$�Rs ���D$8    t����L$ �\$�5s �ƋL$0d�    Y^[��0� ���������������j�h�Ud�    P��8SUVW�  3�P�D$Ld�    �����    �D$u�D$\�t$`��l$`��t$\�l$`��tE�_����	 ��t.�o8����$����t���$���\$����	 �L$�l$`��l$`���D$ ���t]�d tr�L$ �e����Od����   j ���T$,�$R�D$d    �Ѕ�	���D$ �	�L$ �{]���L$ �] �D$T�����G����D$�L$Ld�    Y_^][��D� ��2��] ���ދT$3�8��   ��;�u�   � V�   +�;�^u�yd t�Id��Px��� 3�� VW�|$��t[�T$3�8��   ��;�u'���   j ����"���j���"���__�   ^� �   +�;�u�yd t�Id��P|W��_^� _3�^� ���̋T$3�8��   ��;�uA�D$��t�     �D$��t#���   ����   �P���   �P���   �H�   � V�   +�;�^u/�yd t)�D$�D$�Id����   P�D$P�D$P���$��� 3�� ����������̋T$3�8��   ��;�u�   � V�   +�;�^u�yd t�Id����   ��� 3�� ������������̋T$3�8��   ��;�u�D$�D$P�D$P���$R�#� � V�   +�;�^u*�yd t$�D$�D$�Id����   P�D$P���$��� 3�� ������ �����������U������4  SVW���d �  �Od�E����   ���$�҅��  �u����  �Od��$�   P�l�����$�   Q�Od�ܷ���T$8�_R����	 �GH�OL�WP�D$h�GT�L$l�OX�T$p�W\�D$t�D$8�L$xP�L$l��$�   Q��$�   R�	1������$�   �j0����u��$�   �.��݄$�   �D$hP����$  �$Q��)��݄$�   ��P��$�   R��$�   P����$$  �$Q�)����P��$�   R����(������(��݄$�   �D$hP����$�   �$Q�t)��݄$�   ��P��$,  R��$�   P����$$  �$Q�F)����P��$  R���c(�����\(����$�   P��$�   Q��$0  �p(��P�T$<R�D$XP��/�����L$P�-����$�   ��$�   ��$�   ���$�   �V��$�   �F�N�V��$�   �L$8�T$<�F���    up�D$@�N0�L$D�~0�W�T$H�G�D$L�O��$�   Q�W�L$T�G��*����VH�P�NH�Q�P�Q�P�Q�P�Q�@Q�A��$�   WQ�-/���N�c�F��L$@�P�T$D�H�L$H�P�T$L�H�P�T$P�VH�T$T�NH�Q�T$X�Q�T$\�Q�T$`P�Q�T$hQ��$�   P�Q��.���N0���P�Q�P�Q�P�Q�P�Q�@���A�k,�����$� �   _^[��]� _^3�[��]� �����������3�8��   �   ��+�;T$u�yd t�Id����   ��� 3�� �������������3�8��   �   ��+�;T$u�yd t�Id����   ��� 3�� ������������̋T$3�8��   ��;�uA�D$0�D$$���\$�D$8�$P�D$4�D$(P�D$4P�D$$���\$�D$8�$PR�� �4 V�   +�;�^uN�yd tH�D$0�D$$�Id����   ���\$�D$8�$P�D$4�D$(P�D$4P�D$$���\$�D$8�$P���4 2��4 �����������̃yd u2��@ ���    �D$t�D$����D$t���3��D$<�Id����   ��(�\$ �D$\�\$�D$T�\$�D$L�\$�D$D�$P�D$0���$P���@ ��������������{� ����������́�   V��3�9Fd��   8��   ��$�   ��;�uL���   �m���N�է	 ����$�L$�t����0'�D$�\$j P����������^�Ā   � �   +�;�u�Nd����   ��^�Ā   � 3�^�Ā   � �������������̀��    �����   �   �����������U�������  SV��~d Wu3�_^[��]�$ ���    �E$��   ���E�E�]��   ����   �   �}(�Nd�]����   WP�E P�EPS���$�҅�t��E�����   �$�����T$0�荌$�   ���\$8�������$h  �����D$@�~P���ϥ	 �D$8��$����DzC��?��$�   �n����
  �E���Z������Q�����t��t3��E�������=����~j t	�Np�L$,��D$,    �F8����$�  �$R���l�	 �T$,j j ��$�   QR�VH���̉�VL�Q�VP�Q�VT�Q�VX�Q�V\�Q�T$h���̉��$�   �Q��$�   �Q��$�   �Q��$�   �Q��$�   �Q����̉�P�Q�P�Q�P�Q�P�@�Q�A�Z�����X���&����D$0��$����Dz����$h  �>�����   �~k t���   �L$,��D$,    �F@����$�  �$R���g�	 �T$,j j ��$p  QR�VH���̉�VL�Q�VP�Q�VT�Q�VX�Q�V\�Q�T$h���̉��$�   �Q��$�   �Q��$�   �Q��$�   �Q��$�   �Q����̉�P�Q�P�Q�P�Q�P�@�Q�A�U�����X���!���݄$�   �{���G�D$8����݄$h  ���D$0�������+��\$X�U ݄$�   �����E����݄$p  ����������������\$`݄$   ��݄$�  �������\$h݄$  ��݄$�  �΍<������\$p݄$  ��݄$�  �����\$x݄$   ��݄$�  ����ݜ$�   ݄$(  ��݄$�  ����ݜ$�   ݄$0  ��݄$�  ����ݜ$�   ݄$@  ��݄$�  ��������ݜ$�   ��G����  ݆�   ܦ�   ��������z�����ˋE�����������������݄$�  ܤ$   ��ݜ$�   ݄$�  ܤ$  ��݄$�  ܤ$  ��ݔ$�   ݄$�  ܤ$   ��ݜ$�   ݄$�  ܤ$(  ��ݜ$�   ݄$�  ܤ$0  ��ݜ$�   ݄$�  ܤ$@  ����ݜ$�   �����݄$�   ��������������+��\$0�S������\$8�T$,��Gu��������Q�Q�+ȃ�u��؃�����������u:܄$�   �����������܄$�   �Y݄$�   ��݄$�   ����܄$�   �#������������Y݄$�   ��݄$�   �����Y+��D$8�\$,�L$`�D$0�L$X����D$8�L$x�D$0�L$p���Y�D$8܌$�   �D$0܌$�   ���Y+ȅ�������]�ڋE�����
�����������D$`���D$X�����D$h��D$x���D$p����܄$�   �Y܌$�   ݄$�   ����܄$�   �Y���    ��   ����   ��|�   ��    ���   w��$�   �T$0�S�u������D$0�   9U�   �E����D$,�J�����E�+U ���4D$,�<0;��L$8s8�L$0SVQ�Q�
 SWV�I�
 �T$HSRW�=�
 �E����+���$;�r̋L$8�E���D$,��;U~��D$0��$�   ;�t	P������_^�   [��]�$ �����������U����j�h�Ud�    P��  SVW�  3�P��$�  d�    ��~d u3���$�  d�    Y_^[��]� ���    t�   +E�E�D$�~P��詞	 ��$�   譢���L$4褢���~j t�^p�3��F8����$D  �$Q��菞	 j j ��$�   R�VHS���̉�VL�Q�VP�Q�VT�Q�VX�Q�V\�Q�T$D���̉�T$`�Q�T$d�Q�T$h�Q�T$l�Q�T$p�Q����̉�P�Q�P�Q�P�Q�P�@�Q�A萬����X��������~k t���   �3��F@����$D  �$Q���͝	 j j �T$<R�VHS���̉�VL�Q�VP�Q�VT�Q�VX�Q�V\�Q�T$D���̉�T$`�Q�T$d�Q�T$h�Q�T$l�Q�T$p�Q����̉�P�Q�P�Q�P�Q�P�@�Q�A�ѫ����X���0����E3�����   �E����$\  �$Q�Nd诧��jP�X�������$�   ;ǉ�$�  t	����? �����   ���   �W8�H�O<�P�W@�@��$T  Q��$@  R��$�   Ǆ$�  �����GD�GH   �ۥ����O�P�W�H�O�P�W�H�O�P��$T  P��$p  Q�L$<�W蟥����W �H�O$�P�W(�H�O,�P�W0�@�G4��  ����  �E�����   �$��������݄$�   ���D$4�����\$4݄$�   ���D$<�����\$<݄$�   ���D$D�����\$D݄$�   ���D$L�����\$L݄$�   ���D$T�����\$T݄$�   ���D$\�����\$\݄$�   ���D$d�����\$d݄$�   ���D$l�����\$l݄$�   ���D$t�����\$t݄$  ���D$|�����\$|݄$  ��݄$�   ����ݜ$�   ݄$  ��݄$�   ����ݜ$�   ݄$  ��݄$�   �Nd����ݜ$�   ݄$$  ��݄$�   ����ݜ$�   ݄$,  ��݄$�   ����ݜ$�   ܌$4  ݄$�   ����ݜ$�   ��Bd�Ћ���tO��Btj���Ћ�RD�D$4P���҅�u2��P���$P��觝������Pj���҅���t��PD�L$4Q���ҋǋ�$�  d�    Y_^[��]� ������������U����j�hVd�    P��hSVW�  3�P�D$xd�    �ًu���D$ �c����u3��L$xd�    Y_^[��]� ���    t
�   +E��E����  ���   ��������D$�  V���$������  �L$4����WV�L$<Ǆ$�       �q%���L$4�������D$��  j �L$8���� �����$�����\$j�L$8���� �����$�����\$$�s8j ���d�����d$j����\$ �O��� j �L$���D$ �\$ �8����j�d$(����\$0�#��� �D$$�����D$,�T$$���\$����Aup�D$��$����u]������zV��������uMj ���D$�D$ ����� �D$��������D{0��������z'j ���D$����D$��Cj ������D$ �g��j������ �D$$��������D{ ��������Auj���[���D$$��Ck �	�؀|$ t"�D$4�L$8�T$<��D$@�O�W�ˉG�����L$4Ǆ$�   ������Z �$��u �Kd��t����   V�Ѕ����D$誏���D$�L$xd�    Y_^[��]� U������tSV��M2���W��  �]��������t���   �������u2�_^[��]� j ����������$�����T$ ����������z�\$ ���j���b�������$����T$(����������Au�\$(��؍^8j ��� �����d$ j����\$4���� j �L$$���D$4�\$$��
����j�d$,����\$4��
���D$(�N��F�V�~�D$0�L$<�O�D$8�G�\$(�T$@�W�L$H�N$�D$D�F �T$L�V(�L$T�N0�D$P�F,�T$X�V4�L$`j ���D$# �D$`�T$h�l
��� �\$ ����Au�Mj �D$#�`
��ݞ�   ���D$ ��������zH���D$p�$P���Ǖ	 ��P�L$8�H�T$<�P�L$@�H�T$D�P�L$Hj �ˉT$P��	�����j �؋���	���D$ �j����	��� �\$(����z~�Mj��	��ݞ�   ���D$(��������AuJ���D$p�$P���7�	 ��P�L$P�H�T$T�P�L$X�H�T$\�P�L$`j�ˉT$h�e	������j�؋��T	���D$(���|$ tZ�D$8�L$<�T$@��D$D�O�L$H�W�T$L�G�D$P�O�L$T�F �D$\�N$�L$`�W�T$X�V(�T$d�F,�N0�ΉV4諌���_^[��]� ��u�Nd��t��U���   R�Њ؄�t���z���_^��[��]� ���������������j�hVVd�    P��\  UVW�  3�P��$l  d�    ��}d u3���  �L$l������$�   �������D$lP�����$������t��荌$�   Q�����$������t��L$�I��݄$�  �Md����   j ���D$ �$PǄ$�      �ҋ����t$�L$Ǆ$t  ������w�����)  �|$tj�L$�1F���D$P�L$D�v���L$lQ�L$Ƅ$x  �]L����$�   R�L$D�LL���D$(�L$$�T$ ��$|  jPjQRj����* j ���P� �N(���P�D$4PQ�{�
 �����   j ���9���V,j����+���F,3��X9~~6W�L$��*��Pjj W��� W�L$D�*��PjjW���� ��;~|ʀ��    t����   ���ЍL$@Ƅ$t   �v���L$Ǆ$t  �����v���D$��$l  d�    Y_^]��h  � ��������������̃yd t�Id����   ��3�����������̀��    V�t�D$�t$�D$�T$�\$��t$�D$�T$��t#�yd t�Id�R���   ���$�҅����2��؅�t�D$�^� ����������̀��    V�t�D$�t$�D$�T$�\$��t$�D$�T$��t#�yd t�Id�R���   ���$�҅����2��؅�t�D$�^� �����������j�h�Vd�    P���   SUVW�  3�P��$�   d�    �L$��$�   ��tg�k(�s�   ���t��Pj���    ��=�C��=�K��=�S��=�C��=�K ��=�͉S$�S ����u��L$�yd �  ���L$ �Ǐ	 ���
  �l$���D�������  �L$l�#�����D$lP�����$�O�������  ���D$    蘪������   �MdQ趰 ������tx����'����ulj ���(� ��t_��ȋBd�ЋMd��Rh���D$$P�ҋ���̉�P�Q�P�@�Q�A��Ǆ$      轇���L$$Ǆ$�   �����R ��u�Md��Bd�Ћ����  ���;���   �����$�Ѕ��   W��1 ������   jP�y������D$��Ǆ$�      t����1 ���3��L$$Q��Ǆ$�   ����������V�H�N�P�V�H�N�P�V�@�L$$Q�ωF�`�����V �H�N$�P�V(�H�N,�P�V0�@�F4��Rh�D$$P���ҋ���̉�P�Q�P�@�Q�A��Ǆ$     蒆���L$$Ǆ$�   �����~Q ��Bj���Ћ���Btj���Є���  ����L$t�$�}�����u��RD�D$lP���҅���  jP�L������D$��Ǆ$�      t����0 ���3���Ǆ$�   �����t$�a  ��=�F��=�N��=�V��=�F��=�D$ �N��=P�L$(Q�M �V���P�N ��	���.�L$���   j��l�����L$���$j ���   ����U �����$�҅���   ��uTjX�v������D$��Ǆ$�      t	����E �3��؅�Ǆ$�   ����u��Pj���ҋ�Pj�����   �l$�{�s��=�C��=�K��=�S��=�C��=�K ��=�D$<P�͉S$��� ���{(�   �L$<�O ���    t����   ���Ћ����Bj���ЋL$��t	��Bj��3���$�   d�    Y_^][���   � ������̸K�����������j�h�Vd�    PSVW�  3�P�D$d�    �D$ �����   +��   �> t6h�  �������D$ ���D$    t�Q����j���3��D$�����7����u��L$d�    Y_^[��� ��VW���   �   �I ���t��Pj���    ����u�_^�SV�t$Wh�eV���<� ����貕 ���    ���   u-���    u$���    uh�eV�� ����輕 _^[� 3��d$ �; WuhpeV�ߕ ���&h`eV�ϕ �����E� ���PV�ҋ��t� ������r����b� _^[� ������������SVW���1 �����Ƹ   �   ��    �> t���P�������u��_^[��̋D$VW���   �   �> t
��P�B�Ѓ���u�_^� ���S�\$UV��W�˿   ��W 3��D$�Ÿ   ��t$�|$ t�E �3�P���E ��������r؋�_^][� �������������QSVW���5���3۾   �Ǹ   ��tN�L$�D$P�D$    ��c ����t�L$Q�^�������L$��t�? u��Bj��3�������r�_��^[Y� ������������̋D$h�eP聚 ���   � �����̃��    u!���    u���    u�   3Ʉ������3�3Ʉ����������������S�\$VW�   3����   ��t�> t
���PDS�҃�����r�_^[� ��������j�h1Wd�    PQ�  3�P�D$d�    �L$�L$���D$    t�f�  �L$d�    Y��� ����j�haWd�    PQ�  3�P�D$d�    �L$�L$���D$    t��  �L$d�    Y��� ����j�h�Wd�    PQ�  3�P�D$d�    �L$�L$���D$    t�F�  �L$d�    Y��� ����j�h�Wd�    PQ�  3�P�D$d�    �L$�L$���D$    t�V�  �L$d�    Y��� ����V�t$��th0J���`����t��^�3�^����������������VW�|$��t5h0J���Z`����t%�t$��th0J���B`����tW������_�^�_2�^�������������j�hXd�    PQSVW�  3�P�D$d�    ��t$�A� �N�D$    �4a�˅	 �N8�D$������NH�D$����~p�   ���������y񍎠   �����D$腙���ƋL$d�    Y_^[���V���ȡ���D$t	V�{�������^� ��U����j�hgXd�    P���   SVW�  3�P��$�   d�    �L$L�uH �}3�9_��$   �\$$�\$(�  �G�[��ȃy ��   �y �  �M�[�ыt�X����  ��$�   �H ��P<j j ��$�   Q��Ƅ$  �҅�u�   ��$�   �|$L�}���$�   P�L$P�K �L$(;L$$uh�T$|R��$�   ��	 ��;�D$|����݄$�   ��Az��e������{��������Az!��e����Au�D$(��D$(��������؃D$$��$�   Ƅ$    ��G ��;_������|$$ ��  �D$d���\$�L$<�D$\�$�����D$l���\$�L$L�D$dƄ$  �$����D$$9D$(���$   |�L$,�������t�L$<������ud�L$,�Y�����$����Dz�����Xe�L$<�D$,���\$,�D$4�\$4�'�����$����Dz�����Xe�D$<���\$<�D$D�\$D�L$,�E�������   �L$<�4�������   h�   �������D$(��Ƅ$   thhY���� ���3��D$,j�����j �D$L���X��$  �Y� �D$<j�����j�D$\���X�<� ��}���$��芍����u
��BDW���ЍL$<Ƅ$   �;F �L$,Ƅ$    �*F �L$LǄ$   �����F �Ƌ�$�   d�    Y_^[��]ÍL$<Ƅ$   ��E �L$,Ƅ$    ��E �L$LǄ$   ������E 3���$�   d�    Y_^[��]Ã�DSV�؅�W����u	��_^[��D�U���4  �����  ����  ;~��  �D$\SP���$ ;~�D$�D$�|$��   �D$X��������X   �T$ �ډD$�N�| |d���T;Tu{�D$���tkP���ס  �N�T$�
    �L$X���FËT�PR���2�  ��t:�L$WQj P���Q ��T$ �Ph�X`�D$�D$`����`;F�D$�v�����D$ �T$R�����  �|$ ��   �L$�y3�����   ��$    �T$�J�4���i��   �D$ ����]d�D$$P�<�i��   ����*���P�L$@Q��蝌�����������t@WV����	 ��t3���nI  ��t	�5�XX���ZI  ��t	�5�XX�D$`��t� �T$�D$ �z;��_����D$]_^[��D�]��_^[��D����������U�����E��4S3�;�VW��   ����   �M9Y�\$<��   �A3��9x��   ��H�IdW���$W�i���������   ��Btj����j���K���E��u��3��/��u	���������M���$�?�����u��E�RDP���҅�t!��M���$������u�M��PDQ���ҋE�H�tX�P�|\�ȋD$<����`;A�D$<�1����_^[��]�_^2�[��]��������������U����j�hYd�    P��(  SVW�  3�P��$8  d�    ��}���C  �E���$�2��������*  �E� 3�;�t�M;�  ��RlW�D$8P�����E���L$<�$��$H  �����T$,����������  ��������A��  S�L$8������ �]������  j�L$8������ �]����A��  �E� 3����|$tP������؃����_  �M���tP����������D$�A  ��3�8��   ��9E�/  ��$�   �@}	 ��$�   Ƅ$@  �,}	 �L$TƄ$@  �;����L$dƄ$@  �*����L$tƄ$@  �����L$DƄ$@  �����~8j ��Ƅ$D  �����\$$j������ݔ$�   ����D$4�����L$,�������T$$�$���������  �D$$�D$��������A��  ܜ$�   ������  �D$,����$�   �$�~R���}	 �O��W��$�   �O��$�   �G��$�   ��$�   ��$�   �W��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   �N(��$�   ��$�   ��$�   ��$�   �V ��$�   �F$��$�   �N4��$�   ��$   ��$�   �V,��$�   �F0��$�   j �L$8��$�   ��$�   ��$�   ��$�   �o����E���\$�L$d� �$�7��j�L$8�L���� ���\$�L$t�E�$����D$���\$��$�   �D$4�$����݄$�   ���\$�L$T�D$,�$������$�   ��z	 ���&  ��$�   �({	 ��;����A�	  ��$�   ��z	 ����  ��$�   ��z	 ��;����A��  ��u?h�   �x������D$$��Ƅ$@  tV������Ƅ$@  ���%3�Ƅ$@  ���;ދ�tV�����	��B0j�ЋL$��u3h�   �������D$$��Ƅ$@  tV��菕���D$�3��D$�;�tV跖���	��B0j�Ѝ{�   ��$�   �L$T���   �T$X���   �D$\���   �L$`���   �T$t�S8�D$x�C<�L$|�D$�K@��$�   �SD�x�   ��$�   �L$d���   �T$h���   �L$l���   �T$p���   �L$D�H8�T$H�P<�L$L�H@�T$P�M�PD�U��L$D�Ƅ$@  ��< �L$tƄ$@  ��< �L$dƄ$@  ��< �L$TƄ$@  �< ��$�   Ƅ$@  �< ��$�   Ƅ$@   �< �  �؍L$DƄ$@  �}< �L$tƄ$@  �l< �L$dƄ$@  �[< �L$TƄ$@  �J< ��$�   Ƅ$@  �6< ��$�   Ƅ$@   �"< ��  3�9Fd��  ;މD$�D$,u�Cd��D$�B0j�����;�t�Kd;�t��Bj���Cd    ;�u�Od��B0�L$,j�������t�Od��t��Bj���Gd    �Nd�E����   �D$,P�D$ P���$�҅��[  �T$���5  �D$,���  �Nd;��D$$    t;�t;�t
;�t�L$$���t	��Pj�҅��Fd    u=h�   �A������D$��Ƅ$@  	tV��趒����$@  ���3���$@  ���;�tV���ғ����u7h�   �������D$��Ƅ$@  
tV���i����D$���3��D$���;�tV��苓���D$$�L$�Fd�E�Kd�T$,�M�Wd��9�L$4Ǆ$@  �����h: �   ��$8  d�    Y_^[��]� 9Vdt%��ʋPj�ҋL$,��t9Ndt��Pj����؍L$4Ǆ$@  �����: 3���$8  d�    Y_^[��]� ���j�hHYd�    P��V�  3�P�D$d�    ��t$�� 3���e�D$$���   ���   ���   �D$P�K�M����N�P�V�H�N�P�V� 0�F�0�N�0�V �0�F$�F(   �ƋL$d�    Y^�� ��j�hxYd�    PQV�  3�P�D$d�    ��t$��e�D$    �U������D$�����V �L$d�    Y^�������̋D$����VW��   �$��3��w��   �w�
�   �   S�\$ ��tI�D$P�K�L��P���L���؅�t,hK���N����t;���}����   �9 u����;�|�[_3�^���3��_3�^��Ë���   [_^��ÍI ��y�������S�\$��UVW��}J3�9nt6�~��x��k�h�N��P�U�҃���h;�}�N��PUQ���҉n_�n�n^][� �F;�}m�N��PSQ����3�;FtI�N��+�k�hk�hWR�Q���
 �F��;�}����k�h+�F�P��������h��u�_�^^][� _�V�V^][� ~R���;�|#��+�k�h����N�9�B�j �Ѓ�h��u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� ��������S�\$��UVW��}P3�9nt<�~��x#��i��   �N��P�U�҃����   ;�}�N��PUQ���҉n_�n�n^][� �F;�}y�N��PSQ����3�;FtU�N��+�i��   i��   WR�Q趿
 �F��;�}$����i��   +�F�P���������   ��u�_�^^][� _�V�V^][� ~X���;�|)��+�i��   ����N�9�B�j �Ё��   ��u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� S�\$��UVW��}J3�9nt6�~��x��k�h�N��P�U�҃���h;�}�N��PUQ���҉n_�n�n^][� �F;�}m�N��PSQ����3�;FtI�N��+�k�hk�hWR�Q肾
 �F��;�}����k�h+�F�P���������h��u�_�^^][� _�V�V^][� ~R���;�|#��+�k�h����N�9�B�j �Ѓ�h��u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� ��������S�\$��UVW��}P3�9nt<�~��x#��iۨ   �N��P�U�҃���   ;�}�N��PUQ���҉n_�n�n^][� �F;�}y�N��PSQ����3�;FtU�N��+�iɨ   i��   WR�Q�F�
 �F��;�}$����i��   +�F�P��������Ǩ   ��u�_�^^][� _�V�V^][� ~X���;�|)��+�i��   ����N�9�B�j �Ё�   ��u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� �D$9A}	�D$�.���� �����������j�h�Yd�    PQ�  3�P�D$d�    h�   �|�����D$���D$    t��������L$d�    Y���3��L$d�    Y������������j�h�Yd�    PQVW�  3�P�D$d�    ��h�   �{�����D$���D$    t���W������3����D$����tW���=����ƋL$d�    Y_^�����������̃�(SUV�t$8Wh<gV����y �����^y h4gV��y ���_8j �ˍo�1������D$(�$P���n	 P���| h0gV�y ��j��� ������L$(�$Q���~n	 P���V| h�&V�ky h(gV�`y ���WHR���} h�&V�Gy �Gi�OhPQhgV�2y �Wk�GjRPh�fV�y h�fV�y ��0�OpQ����| h�fV��x �����   R���| h�&V��x �����   j���;������$j ���,������$h�fV�x ���   Ph�fV�x �O`Qh�fV�x h�fV�~x ��8����w �d uh�fV�cx ����Od��BV�Ћ��x 3��D$   �D$   �D$   �D$ �f�D$$pf�D$(`f�\$��    �LQW�U��������to���D$<Xf轹���؅�t2h A���+�����u
�D$<Pf�h�A��������u�D$<Hf��� �T$�L$<P�D$PQh,fV�w �\$$�������\$�m������6w _^][��(� ������������j�hZd�    PQ�  3�P�D$d�    h�   �x�����D$���D$    t���[����L$d�    Y���3��L$d�    Y������������j�h;Zd�    PQVW�  3�P�D$d�    ��h�   �x�����D$���D$    t����������3����D$����t;�t���
���W���� W���j����ƋL$d�    Y_^���������VW�|$��tHhK���D����t8�t$��t0hK���rD����t ;�t������W���[ W������_�^�_2�^����������V��������D$t	V�;y������^� �̋D$9A}	�D$������ ����������̋D$9A}	�D$������ ����������̋D$9A}	�D$����� ����������̋D$9A}	�D$����� �����������SUVW�|$����}S3�9n�
  �~��x"������    �N�趷������`;�}�N��PUQ����_�n�n�n^][� �F;�}j�N��PWQ����3�;ŉF��   �V��+ʍI�R��Q���UR�O�
 �F��;�}�@����+�N�t蟷����`��u�~_^][� ~U���;�|&�@+������荤$    �N��������`��u�9~~�~�N��PWQ�Ή~��3�;ŉFu�n�n_^][� ���������������QS�ًCd��W�{du_3�[Y� �K`��|�UVu*�t$�F��9F}P������W���V���C`^]_[Y� P草 �����D$tc�s`��� ��;�uU�|$�o�V������3�9s`~��L$V�� ���D$t�D$P���>V����;s`|ڋC`^]_[Y� ��|;o�o^]_3�[Y� ����̋D$V��3�;��Pg�N�N�N~P���������^� �����̋Q2���t%�I��~V�t$��t��~Vj`QR��% ���^� ��������������̋Q2���t%�I��~V�t$��t��~Vj`QR�x% ���^� ��������������̋D$�L$�@��PQ�[������ �����UW��3�9o�Pgt7V�w��xS�v���O���������`;�}�[�O��PUQ���҉o^�o�o_]����������������V�������D$t	V�[u������^� ��V��F�V�@��;�uJ��   v��|�]U ;�}�������   ��;�}7P���W����N�I��F���N^�N�+����F�@��Nt舴���N�I��F���N^�����U����j�h�Zd�    P��h  SVW�  3�P��$x  d�    �ًM3�;�t�n�  �,%�t$d�|$h�|$l�|$p�D$dP�ˉ�$�  ��������D$H��  ;D$l��  ��$�   �sQ���e	 ��$�   �a�����u5h�hh�hh7
  h�e�� ���L$dǄ$�  ����������  �����$L  �$��i������$��$�  �i������$��$L  �i������$��$L  �i������$��$�  �ti������$��$�  �`i���{j t�{p�C8����$�   �$R����d	 ��$�  Q��$H  R�SH��$L  QW���̉�SL�Q�SP�Q�ST�Q�SX�Q�S\�Q��$�   ���̉��$�   �Q��$�   �Q��$   �Q��$  �Q��$  �Q����̉�P�Q�P�Q�P�Q�P�@�Q�A��r����X��uh�hh�hh>
  �y����{k t���   �3��C@����$�   �$Q���d	 ��$�  R��$H  Q��$�  R�SHW���̉�SL�Q�SP�Q�ST�Q�SX�Q�S\�Q��$�   ���̉��$�   �Q��$�   �Q��$   �Q��$  �Q��$  �Q����̉�P�Q�P�Q�P�Q�P�@�Q�A��q����X��uh�hh�hhD
  �����u��t�t$<��u0 ���D$<��uh`hh�hhL
  �Y�������x�����D$4|	����  3��D$43Ʌ����L$8�T$8�D$H�<�N0W��� ���   W�N����|$8�W�T$H�NpR�������|$H�NW�� �N`W������|$H��W�N �� W�NP�������    �   �   ��$�   ��$�   Ǆ$�       ��$�   Ǆ$�      ��$�   t9���   ��$�   ��$�   ��$�   Ǆ$�      ��$�   Ǆ$�       �|$H�?P�L$x������Ƅ$�  �D$@    ��  �L$h�T$@�<�����  �D$|��$�   �D$L路����$�   Ƅ$�  裯����Bd���Ћ����	  ����   ���Ѕ�������$�   t j V��   ����h����D$8   �f���3�3�9L$4��$�   t3�9L$@�T�;�t�L$4�L$8�} ��  �5��$�   Pݔ$�   ��$�   ݜ$�   Q���uX������  ݄$�   ���$�����������  ݄$�   ���$�����������  ݄$�   ݄$�   �������g  �ɋݔ$�   ��4���   ���\$��$�   ��A���$j j P���\$�$j�҄���   ݄$�   ܔ$�   ����A��   ݄$�   ������A��   3��L$`Q��$�   ��$�   �D$d����   R�����$�ЋL$`����$�   tW��tf��tO�L$t�������$�   �HǄ$�       ��Bj����݄$�   �t$`ݔ$�   ݄$�   �D$`    �������t��ȋBj�ЋL$`��t��Bj����؍L$t�a����L$L�p�D$|;ȉD$\�F  ���@���L$P��$�   ��$    �L$x��$�   �
h�   �D$X�@�����]k�����D$X��Ƅ$�  t	�������3��T$T�B�x�   �s�B�K8�H8�K<�H<�K@�H@�KD�HD�KH��8�B�HH�KL�HL�KP�HP�KT�HT�KX�HX�K\�H\��H�B�@`   �J�B�Ad�J�Ah �B�@i �Cj�J�Aj�Ck�J�Ak�B�Kp�Hp�Kt�Ht�Kx�Hx�K|�H|���   ��p�H���   �H�B���   ���   ���   ���   ���   �   �H���   �H���   �H���   �H�B���   �   ����   �H���   Ƅ$�  �H���   �H���   �B��$�   ���   ��$�   �D$@�B��$�   �
��$�   �B����   ��$  �B��$�   �z�L����  ����$�   �D�(|3�9��  ���D�8��$�    t^�D$P;D$L~T�L$\���;�uI��$�   ��$�   �D���$�   ����   �J ��$�   ���  ���D�(|3�9��  ���D�8��t$T�Nj j ���$j �׃ ���D$T��  �N8Q�L$@�V(RWP��	 ���D$Xu�L$T��Bj���T  �L$X�D$P;D$L�Q�Vu8��$�   ��T���$�   ����   ��$�   �L�(�T�8���  ���  �|$4 ��$�   �L��V ����   ��$�   �L�(��$  �T�8���  ���  ��   �|$X���'  ����   ���'  ������   ����$  ����   ��$�   P���Js  3�;��D$Xtb�xPu\��$�   Q���+s  ����tQ�PuK�L$X�$  �ωD$T��#  �|$T t0��t,�T$X�J8�NH�W8�L$T�VL�Q8�VP�@8�FT��L$4�L$8�
3��D$4�D$8�D$P��$�   `��;D$\�D$P�������$�   Ƅ$�  艨���D$@��;D$H�D$@�����t$<�|$4 �D$G ��  3Ƀ|$4����9L$8��  �L$4��$D  R��$H  PQ��$�   R����������  �F8�|$8�P�N0�� ���   �P���   �����3��|$4�D$P�D$Lt�|$4u<��$�  P�L$xj Q��������t!P���+{  P�����  ���    �D$P�P0�D$4��t��u<��$�  P�L$xjQ���������t!P����z  P���y�  ���    �D$L�P0�|$P u�|$L ��  �|$8�L$|�F���Q�N�� �Fx���T$H�R�Np������L$|�Fh���Q�N`�����D$@    �L$@�ɋD$Pt�D$L���D$\tq3�3�9|$H~O;t$|}M�D$x�v��9|u9�T$@3������L$GQ�΃�P�D$dR��$�   ������;�~��;|$H��|�;t$|�p  ;|$H�f  �L$@�����L$@�k����  hHhh�hhx
  h�e�� �L$L��;Mt	��Bj�ЍL$tƄ$�   ���������h hh�hh�
  h�e�`� ���L$<;Mt	��Bj�Ѝ�$�   Ƅ$�  �ץ���L$tƄ$�   ������������hhh�hh�
  h�e�� ��B��j�����h�gh�hh�
  h�e�ۿ �L$L��;Mt	��Bj�Ѝ�$�   Ƅ$�  �R����L$tƄ$�   �1����|$p Ǆ$�  �����D$d,%��  �D$h����  j �p  h�gh�hh�  h�e�W� �D$`�t$L����t
j P���c  �D$L��t
j P���c  ���% �L$@��u'9L$8u!�|$4u�t$<3�8��   �������   ��t$<���    ~h�~X~bS��蚣����Ppj���Ҁ|$G t	j���_  �L$tƄ$�   �>����L$dǄ$�  �����
����Ƌ�$x  d�    Y_^[��]� h�gh�hh�  h�e�g� ��;u�$�����Pj���ҍL$tƄ$�   ���������h`gh�hh.
  h�e�!� ��9|$pǄ$�  �����t$dt�D$h;�tWP�L$l�8%3���$x  d�    Y_^[��]� ����������̋D$jP�d���� �V�t$��thL����.����t��^�3�^���������������̸L�����������VW�|$��;�t-W��0 �G �F �O$�F,�@�N$�W(�N,�V(�W,R���G@�^@_��^� VW�|$��F(Ph|iW�9` ����V���c h�&W� ` ��_^� �������̋D$�Q��Q�P�Q�P�Q�P�Q�I�P�H� ������V�t$��th M���.����t��^�3�^���������������̸ M����������̸   �����������VW�|$��;�t?W� �G0�F0�O4�N4�W8�V8�G<�F<�O@�FH�@�N@�WD�NH�VD�WHR���GX�^X_��^� ��������������SVW�|$W��� ���Ä�u����   h�jW�_ ��_^��[� �F8��}"����   PhPjW��^ ��_2�^��[� �F<��}��t|Ph$jW�^ ��_2�^��[� �F@��}��tWPh�iW�^ ��_2�^��[� �FD��}��t2Ph�iW�o^ ��_2�^��[� �~` u��th�iW�L^ ��2�_^��[� �������������̋A8�L$Ph�jQ�^ ��� �������V�t$��th�M���;,����t��^�3�^���������������̸�M������������ ��   ������SV�t$��;���   WV�� �F0�C0�N4�K4�V8�S8�F<�C<�N@�K@�VD�SD�FH�CH�NL�KL�VP�SP�FT�CT�NX�Cp�@�KX�F`�[`�Kp�Fh�[h݆�   ݛ�   ݆�   ݛ�   ���   ���   �VpR�Ёƀ   ���   �   �_^��[� �������������V��~8 }"�D$��th8lP��\ ���ܷ ��^� �F<��}#�L$��tPhlQ�\ ��買 ��^� W�|$W� ��u����   h�k�   �F@��}�~Pt����   Ph�k�p�FD��}��tnPh�k�]�FH��}��t[Ph�k�J�FP��r��tGPh`k�6��u��t6Phk�%�FT��r��t"Ph�j��FX��} ��tPh�jW��[ ���� _��^� ���    u��th�jW��[ ���Ƕ _��^� _�   ^� ����̋A8�L$PhPlQ�[ ��� �������V�t$��th�N���)����t��^�3�^���������������̸�N�����������SV�t$��;�tBWV�M4���F�C�N�C�@�K�V�K�S�VR�ЋN$�K$�V(��0�{0�   �S(�_^��[� ����������̅�tQhdlP��Z ���������������V�t$��th�O����(����t��^�3�^���������������̸�O�����������j�h�Zd�    PSVW�  3�P�D$d�    ��|$ ;��a  W��+ �G�F�O�F�@�N�W�N�V�WR�ЋO,�N,�W0�V0�G4�F4�O8�N8�W<�V<�G@�F@�OD�ND���   3�;�t��Bj�Љ��   9��   t9h�  �1[�����D$ ;É\$t���   Q����-���3��D$�������   ���   ;�t��Bj�Љ��   9��   t=h�  ��Z�����D$ ;��D$   t���   Q���-���3��D$�������   ���   ;�t��Bj�Љ��   9��   t5h�  �yZ�����D$ ;��D$   t���   Q���(-���3����   �ƋL$d�    Y_^[��� ������̋��   ����������V�t$W���GPh�lV�X ��8h`/W�q������t$h�lV�X ��W����^ h�lV�X ��h�&V�uX ��_^� ������������̊T$�D$V����I ��ts��tI��tjj�������jj���������   �ҋ��   ��ta��t	��Pj��ǆ�       ^� ���   ��t<��t	��Pj��ǆ�       ^� ���   ��t��t	��Pj��ǆ�       ^� ��̸�P�����������j�h[d�    P��xUVW�  3�P��$�   d�    ��$�   �L$(��������   �   �|$X�Ǆ$�       �D$p�����D$X��������4����;������Au�����������\$X�������\$p�D$x�����D$`������������������z������ʍD$��P���\$d���\$|��V����L$(�P�T$,�H�L$0�P�T$4�H�L$8�Pj �D$,P�L$`�T$D�� ��u1��t�M8QhmS�yV ���L$XǄ$�   ����� 2��H  �T$R����V����L$(�P�T$,�H�L$0�P�T$4�H�L$8�Pj �D$,P�L$`�T$D�F ��u1��t�M8Qh�lS��U ���L$XǄ$�   ����� 2���   �U �Rh�D$P������$�����$Ƅ$�   �7������D$H�$P���EU����L$(�P�T$,�H�L$0�P�T$4�H�L$8�P�L$�T$<Ƅ$�    � j �D$,P�L$`� ��u.��t�M8Qh�lS�DU ���L$XǄ$�   �����] 2���L$XǄ$�   �����E ���$�   d�    Y_^]�Ą   ����������̋D$����ǁ�       w5�$���ǁ�      �"ǁ�      �ǁ�      �
ǁ�      �|$ t
���   � ���   � ��=�I�U�a��������̸   ����������́��   � ����̃�H� ��������U����j�h\[d�    P��(  SVW�  3�P��$8  d�    ��$�   �RN 3���$�   ��$@  �=����$�   ݜ$�   Ƅ$@  �`����L$T�W����E;��A  ��u;���2  V�gi �؃�;߉�$�   �[  ���|������L$t�t$p�ͼ����$�   Ƅ$@  蹼����Ƅ$@  �|$P��  �u��W��$�   P��谆 ��L$t�P�T$x�H�L$|�P��$�   ��$�   �F j�L$x�k���j �ΉD$H�n����D$D������  j �L$x�B���j�ΉD$H�E����L$D�����A��  W���� ����Rh��$�   P���ҋ��$�   �P��$�   �H��$�   �P��$�   ��$�   �
 j �L$x�˻��j �΋��л�������At#j�L$x謻��j�΋�豻��������  j �L$x艻��j �΋�莻���j ����Au	���|�����L$x�a���� j�\$H�L$x�P���j�΋��U����j����z	���C�����L$x�(���� �D$tݜ$�   P��$�   �>�����ti�D$D���L$|�$�W����\$D݄$�   ���L$|�$�=���ݜ$�   �D$D����$�   �$�����\$D݄$�   ����$�   �$�ú���݄$�   ���\$��$�   �D$T�$�`����U��$�   Q�MR��$�   PWQ���������tT�E� �|$P܄$�   ��$�   ���;|$p�|$P�������$�   Ƅ$@  �� �L$tƄ$@  �� ��  ��U��$�   �Ƅ$@  � �L$tƄ$@  � ��$�   Ƅ$@   � ��$�   Ǆ$@  �����pL 3���$8  d�    Y_^[��]Ë�Px���ҋ؃��\$p|�����   ���ҋ����|$D
�D$D   �6��}5��    ���D$D   }���$    ��L$D�	�D$D�Ã�|�|$D�TR��$�   �K ����\��   ;��\���$�   �D$P~�D$D�D$P��;ǉD$P���\��|��؋�P|Q���҅�������}���EtP��$�   Q���M����T$T�H�L$X�P�T$\�H�L$`�P�T$d�@�D$h3�9D$p�D$P�J  �
��    �D$P��$�   �D����\$����$�   �$�(���j��$�   �:����Mj ���>����������  j ��$�   �����Mj�����������A��  j��$�   �����Mj�����������z�Mj�ݷ��ݜ$�   j ��$�   踷���Mj ��輷�������Au�Mj 詷��ݜ$�   j ��$�   脷��j��$�   ���t���� �����A�  3�9t$D�  ���$    �L$T�T$X�D$\��$�   �L$`��$�   �T$d��$�   �D$h��$�   ��$�   ��$�   �����$�   �$��������$�   �$Q�M�#M������T$T�H�L$X�P�T$\�H�L$`�P�T$d�@�D$ht=�L$TQ��$�   R���K����L$T�P�T$X�H�L$\�P�T$`�H�L$d�P�T$h�D$\��;t$D܄$�   ݄$�   �d$T��܄$�   ݜ$�   ������D$P��;D$p�D$P������u�L$X�D$T�T$\��$�   �L$d��$�   �D$`��$�   �T$h��$�   �Mj��$�   ��$�   ��������$�   �$P���L������L$T�P�T$X�p�t$\�X�\$`�X�\$d�@�D$h�E��L$`�P�T$h�p�H�X�Pt=�D$TP��$�   Q���PJ����T$T�H�L$X�P�T$\�H�L$`�P�T$d�@�D$h�D$\�M܄$�   ݄$�   �d$T��܄$�   ݔ$�   ��$���$�   Ƅ$@   �� ��$�   Ǆ$@  �����G �   ��$8  d�    Y_^[��]�j�h�[d�    P��0SVW�  3�P�D$@d�    ��t$P�D$(�\$P��3���K����Rh�D$P���ҋ|$T;��\$Ht������$�iJ����t3��D$PW�L$ Q�T$4VR��������t&���D$������Au�ػ   ���������z����L$�D$H������ �ËL$@d�    Y_^[��<��������������������������� ����������̋D$VP������NH� ^� ������̸   �����������U����j�h�[d�    P��8SVW�  3�P�D$Hd�    ��~0��������؄ۈ\$��   �L$� �} �D$P    tT�u��]�\$W�F�L$�\$ ���T$(��\$0�C�\$8�\$@�/ �D$��D$�^�D$,��D$4�[�\$���E��F8�X�E�FH��FP�X�L$�D$P����� �ËL$Hd�    Y_^[��]� ����������̋A(V�t$Pj���m	 ��^� �������̋A8V�t$Pj���m	 ��^� �������̋AV�t$Pj���nm	 ��^� �������̋A8V�t$Pj���Nm	 ��^� �������̋AV�t$Pj���.m	 ��^� ��������V��F��t�N��Qj P��
 ���F    ^����������̋D$VW��3�9~~S3ۋN��P�B�Ѓ���H;~|�[_^� ��������������̋D$VW��3�9~~S3ۋN��P�B�Ѓ���h;~|�[_^� ��������������̋D$VW��3�9~~ S3ۋN��P�B�Ѓ��è   ;~|�[_^� �����������̋T$V�t$�W�:��+�x���B+Fx���B+Fy_���^�+�x���F+Bx���N+Jy_�   ^�_3�^�����̋Q2���t%�I��~V�t$��t��~VjHQR��� ���^� ��������������̋Q2���t%�I��~V�t$��t��~VjHQR�� ���^� ��������������̋D$�L$�����PQ�b����� �̋Q2���t%�I��~V�t$��t��~VjhQR�H� ���^� ��������������̋D$�L$k�hPQ�.b����� �������̋Q2���t%�I��~V�t$��t��~VjhQR��� ���^� ��������������̋Q2���t(�I��~!V�t$��t��~Vh�   QR�� ���^� �����������̋Q2���t(�I��~!V�t$��t��~Vh�   QR�e� ���^� �����������̋D$�L$i��   PQ�Ka����� �����VW�|$��t5hL�������t%�t$��thL�������tW������_�^�_2�^�������������V���h���N8��@��^��������������VW�|$��t5h M���*����t%�t$��th M�������tW���6���_�^�_2�^�������������V���h� �FT��8   ^�������������j�h\d�    P��xSVW�  3�P��$�   d�    ��3ۉ\$� ���D$uz�F@��|s;FDun���& ��tc���& ��Rh�L$0Q���ҋ���$�   �D$ �   P�Ή\$��� ��$�   �   W�ȉ\$�������t�F`��t�@H9F@�D$|�D$ ��Ǆ$�       t����L$ �\$��� ��Ǆ$�   ����t	�L$0��� �|$ ��   �F@�N`���AD�L$XQ�΍<��C���T$pR���D���G�D$@�O�L$D�W�T$H�G�D$L�O�L$P�W�T$T�G@�D$p�\$P�L$\�I����^X����Az7�L$XQ�L$D�1����\$����Az�T$pR�L$D�����\$����A�   {�D$��$�   d�    Y_^[�Ą   ������������VW�|$��t5h�M��������t%�t$��th�M��������tW�������_�^�_2�^������������̋��   3���t�I@��|;JX}k�hJT������������������VW�|$��t5h�N���j����t%�t$��th�N���R����tW������_�^�_2�^�������������V���8���N ��`��^�������������̋A�������������V��N��}.�t$��tQhdlV�A hDnV�A ��菜 ��^� �   9F}�t$��t�QhdlV�jA h,n��W�~$��wd�~( }.�|$���Y�����tr�F(PhnW�6A ���.� _��^� �~` uU�t$���%�����t>h�mV�A ����� _��^� �t$��tQhdlV��@ Wh�mV��@ ���Λ ��_^� �����̋A�Q$P�A(�IR�T$PQh\nR�@ ��� �����������VW�|$��t5h�O�������t%�t$��th�O�������tW�������_�^�_2�^�������������VW���W �N(�   ���    �<�t���   ��B������    t���   ��B������    t���   ��B�����_^���������������̋A$�������������S�Y$UV3���W~-�y ���|���   ;Bx}�Rt��k�h�|*$t����;�|�_^]3�[Ë��   k�hAt_^][��������������̋A��}�L$��tPh,oQ�E? ��3�� �y$}�D$��th�nP�$? ��3�� �A,��}�L$��t�Ph�nQ�? ��3�� ���    u�D$��t�h�nP��> ��3�� �   � �������������V�t$��th�P��������t��^�3�^����������������QSUVW�������N<N,�^N�   ��3��ۉT$~"��    �F����t��B��D$��;�|�^(3���~�N$����t��B��D$��;�|�^83���~"��    �N4����t��B��D$��;�|�nH3ۅ�~3��ND�9�B���؃�H��u�FL+FH���FX��T$3ۅ�~!3�����I �FT���B��؃�h��u�N\+NX�nhk�h�L$3ۅ�~3��Vd���P��؁��   ��u�Fl+Fh�nxi��   �D$3ۅ�~3���    �Nt�9�B���؃�h��u�N|+Nx���   k�h�L$3ۅ�~ 3����   ���P��؁Ǩ   ��u⋆�   +��   _i��   ^�D$][Y�V��L$�F(PjQ譖 �V@RjP衖 �V4�N0�Q�RP菖 ��$^� �������̋D$VP���S� �N8QjP�g� �V<RjP�[� �N@QjP�O� �NP�VL�R�QP�=� ��XVjP�1� ��<^� ���������̋D$VP���S �NQjP�� �V0RjP��� �V$�N �Q�RP�� ��$^� �̋D$V��P�N@�p���P�NP����P���   �����^� �������S��W���   ��~2U�l$V3����$    ��D$���   PU��-����ƨ   ��u�^]_[� �����������3�9AH��������j�hH\d�    P��SUV�  3�P�D$d�    ��F4�\$,�,��L$����D$(6U�L$�D$(    ��� j W�L$��� �N4�<����   �����   ~F�D$��I �\$,9^,t���0 ;�u���� W�Ί�� ��t���p �ƨ   �l$uÅ�t�U �Bj���ЍL$�D$$�����2���L$d�    Y^][������������������V��~ �dot%�F��tj P�po�F    �F    �F    ^�����������VW�|$��;�t?�G��_�F    ��^� 9F}P�4���N��t�G�F�W��PRQ�x
 ��_��^� ��������������V��~ �Tmt%�F��tj P�`m�F    �F    �F    ^����������̃|$ V�t$t:�FP����   U�nX����   ;ix��   ��k�hQt�R$��u]�   ^� 3��̓�u]�B^� �V@���u]�B^� ����   ;QX}}k�hQTSW�zP��u�ZL�;^8u	��_[]^� ��~S�   3ۅ��D$~D�F8�rL�D$�;T$t��|;Qh}�Adi��   9lXt�D$����;�|�_[]^� �   _[]^� ����������j�h�\d�    P��4SUVW�  3�P�D$Hd�    �ًl$X���  ;kh�  �t$\��i��   {d9o8t=���  UhzV�8 �����7 �G8UPh�yV� 8 �����7 ��  ��BV���Ѕ�u����  UhzV��7 ���  �G<���P  ;C�G  �K�����D$u-����  UhzV�7 �����7 �<WWh�y�r����ȋ�B4�Ѓ��D$\tB���H  UhzV�R7 ������6 �L$\�<QWWhhyV�37 ������6 �  ���} 9D$t8����  UhzV�7 �����y6 h<yV��6 �����6 ��  ��Rh�D$(P���ҋL$��@h�T$8R�D$T    �ЍL$(�D$P�+�������   ��tQUhzV�6 �����	6 j�L$,�ޟ��j �L$,���џ������\$� �$h�xV�X6 �����6 �I� �L$8���D$P �i� �L$(�D$P�����X� ���  j �L$,Q�L$@豢������   ��t�UhzV��5 �����o5 j�L$<�D���j �L$<���7���j�L$,���*���j �L$,�D$\������W<�L$X���\$�E �$R����\$� �$h�xV�5 ��,�.����OD�ɋWH�L$�T$\��
  �CH;���
  ���x
  ;��p
  �GP���W@�T$�D$ ������   ���t6�������UhzV�5 �����4 �T$Rh`xV�5 ������;L$\t;�������UhzV��4 �����X4 �D$\�L$PQhxV��4 ���f����L$����   �Ѕ���  ���O����L$XQhzV�4 �����4 �<WWh�wV�s4 ���������F  ����  ;CX��  ��GLk�hkT3҄���9L�@t:��������T$XRhzV�4 �����3 �D$PhxwV�4 �������T$\3Ʉ���9T�@t:��������D$XPhzV��3 �����J3 �L$Qh8wV�3 ���]����T$8R�L$,蔳����t_�L$����   �҅�tM�D$\9D$tC���.����L$XQhzV�l3 ������2 �W<�D$\�L$RPQh�vV�I3 ��������UP3���~#�ML�l$X�L$\9)t����;�|�����D$ }:��������\$XShzV��2 �����s2 �W@RSh�vV��2 ����������   �D$\3�9(��������   ;Ch��   ;���   i��   Cd�PX;WXu~�Ptx���>�����PhzV�~2 ������1 �OX�W@QRhXvV�a2 �������������D$XPhzV�A2 �����1 �[X�O@SQh�uV�$2 ��������GX����  ;Cx��  �O@��|@�|$  }9��������T$XRhzV��1 �����X1 �G@Ph�uV��1 ���l����WP���a  ���$�%�����T����L$XQhzV�1 �����1 hhuV�}1 ��� ���k�hk�hKTCt�yP~;���������T$XRhzV�I1 �����0 �G@Ph uV�01 ��������@$���  ���  ����������L$XQhzV��0 �����o0 �WXRh�tV��0 ������k�hk�hKTCt�yP};�����n����D$XPhzV�0 �����"0 �O@QhxtV�0 ���6����@$���{  ���r  ���������T$XRhzV�\0 ������/ �GXPh(tV�C0 ���������k�hSt�T$$��k�hST�T$�RP���T$};����������L$XQhzV��/ �����s/ �W@Rh�sV��/ ������3���D$�����l$\~o9l$ tO�T$�RL�,�;l$X��   ���  ;kh��   ��i��   Sd�zPu9BXu�T$����   �l$�l$\�T$��;�l$\|��|$ ��   ���������L$XQhzV�A/ �����. h�sV�,/ ����������������Qh�sV�/ �����. �D$X�L$\�T$ PQRhtsV��. ����������������D$XURPhHsV��. �����<. �OX�W@QRhsV�. ���L��������I���Qh�sV�. �����. �D$\UPh�rV�p. �������D$$�x$�V  ���M  ����������L$XQhzV�7. �����- �WXRh�rV�. ��������GT���  ����   ����   ����   ����������D$XPhzV��- �����K- hHrV��- ���c���k�hCt�x$u�G<��|;C}��|	;KX��   ���>���k�hCt�x$u���u�9O<u�݇�   ܟ�   ����Dz�݇�   ܟ�   ����Dz�݇�   ܟ�   ����Dz��5ܗ�   ����D�[  ܟ�   ����D�L  ܗ�   ����D�;  �W`����Au@����������L$XQhzV��, �����V, �G`���$hrV��, ���e����_h����Au>���Z����T$XRhzV�, �����, �Gh���$h�qV�z, ���������   �W�����u5�������D$XPhzV�K, ������+ h�qV�6, �������9��   t5��������L$XQhzV�, �����+ h�qV��+ �������L$8�D$P �� �L$(�D$P������ ��  �����t��������j����T$XRhzV�+ �����+ hHqV�+ ���6��������3����D$XPhzV�q+ ������* h�pV�\+ ���������������L$XQhzV�<+ �����* h�pV�'+ ���������������T$XRhzV�+ �����}* �[x�GXSPhdpV��* �������������UhzV��* �����D* �[H�L$\SQUh$pV�* ���R������Q���UhzV�* �����	* �[H�T$SRUh�oV�t* ��������tRUhzV�\* ������) �C�O<Pj Qh�oV�=* ������) ��D$\��t�ShRUhxoP�* ���� �L$Hd�    Y_^][��@� �I d�8�� X!�!N#�#����U����j�h�\d�    P���   SVW�  3�P��$�   d�    �ى\$D�u����  ;sx��  ��k�h{t9w�|$Pt@�]����  VhdlS�\) ������( �GVPh�}S�B) ������( �O  �G(����  ;��   ��  �O�ɉL$L;�}���"  VhdlW��( �����p( h`}W��( �����( ��  �G$��tO��tJ��tE�]����  VhdlS�( �����#( �O$jjjQh$}S�( �����D( �  9_`t+�}����  Vh }W�c( ������' h�|�d���3���~c�G��3ۅ��L$H~9�(  ����;�|�]SQ�L$L�������M  �T$H�D$Di��   �Hd�E9D
X�`  ��;t$L|��\$D�$ud�G���5  �Ё�  �yJ���B�   3Ʌ�~=�Sd�G�I �0�t$Ti��   �~P�[  �vT��|	����  ����;O|̍L$|������$�   �����3�9D$L�D$H�  �O0�?�������  �u���X  �EPhdlV�-' �����& h�|V�' ������& �%  �}���  �URhdlW��& �����e& �D$HPSVhp|W��& �����& ��  ����  �MQhdlS�& �����#& �T$HRVhD|�K�������  PhdlS�& ������% �E�T$D�RdP�D$L��i��   �LXQPVh|S�L& �����& �Y  �}���L$H�J  �EPh�{W�& �����% �NP�T$T�D$HjQRPh�{W��% �����% �  �u���L$H��  �MQh�{V��% �����C% �T$T�D$HRPhX{V�% �����d% �  �u����  �MQhdlV�% ������$ �WRh({V�l% �����"% �y  �D$H�\$D�O�4���i��   �D$T��|$L�[d��<�i��   �L$l�T$X�PhQ����ҋ�Ph�L$\Q��Ǆ$      �ҋD$D�@�v<�<�4��<�j�L$pƄ$  �;���� ����$�   �$Q���d$����T$|�H��$�   �P��$�   �H��$�   �P��$�   �@j �L$`��$�   ����� ����$�   �$Q���
$����;���$�   �H��$�   �P��$�   �H��$�   �P��$�   �@��$�   ���$��$�   Q��$�   R��$�   藖����� �������   ݄$�   �����D$|������� {��݄$�   ����݄$�   ������������;������Au������������Au�������������������������������AtI������AtD�L$\Ƅ$    �� �L$lǄ$   ������ �D$T;D$L�|$P�D$H�������������؋u����   �EPhdlV�# �����" ݄$�   �|$P�D$H�O�����\$݄$�   �$RPh�zV��" ݄$�   �D$x�\$�O݄$�   ���\$��RPh�zV�" �� ���`" �} �L$\��Ƅ$    �� �L$lǄ$   ������ �Ë�$�   d�    Y_^[��]� ���$�   d�    Y_^[��]� �u��tU�MQhdlV�*" �����! ���   �G(RPhpzV�
" ������! ��E��t�KxQVh0zP��! ����| ��$�   d�    Y_^[��]� ������̃�U�l$��L$��  ;��   ��  S��iۨ   ��   V9k�t$ �\$tF����   Uh|�V�o! ������  �CUPhT�V�U! �����! �F| ^[]��� 9��   t!��tWUh|�V�%! �����  h(��*�C$���D$=��t+Uh|�V��  �����o  h�V��  �����  ��{ ^[]��� W3�����   ��C ��3��~�d$ 9�   ����;�|�L$VS��������  �L$��k�hit9]�=  �D$ 9E(�g  ��uE�}$tP��t,Ph|�V�O  ������ Sh�V�9  ������ �*{ _^[]��� �m$��t	���J  �\$��;|$�>�����{,����  �D$;x8��  �H4�<� ���D$ �>  ��t�Uh|�V�� �����6 �S,Rh��i������q����T$ Rh|�V� ����� SUWhXV�x ���:������9����D$ Ph|�V�X ������ SWh(V�A �������������L$ Qh|�V�! ����� SWhV�
 ��������������Ph|�V�� �����d �T$ �E(RPSSWh�~V�� �������������Ph|�V� �����' SWh�~V� ���\�������  �L$ 9t)���L���Uh|�V�o ������ WhX~�������#� ��t1������Uh|�V�; ����� h,~V�& �������_^[�]��� �������Uh|�V�� �����t �T$�B8�K,PQh�}V�� �������D$��t���   RUh�}P� ���x ]��� �����������j�h�\d�    P��8SUVW�  3�P�D$Ld�    ���|$(�l$\����  ;oX�x  �t$`��k�h_T9{`�\$t8���v  Uh(�V�5 ����� h��V�  ������ �F  9k8t=���9  Uh(�V�� �����n �C8UPhԃV�� ����� �  ��BV���Ѕ�u(����  Uh(�V� �����# h���s����C<���o  ;G(�f  ��    �G$��L$ �ˉD$`��� �L$`9�  �W$�D$ �< ��  �L$,Q�T$8R���������   ���a  �D$<P����� Uh(�V�D$`    � ����� j�L$@�W���j �L$@���J�������\$� �$h��V�� ����� �L$<�D$T������� ��  �C@���SD�K@�D$ �T$`��  �WH;���  �D$`����  ;���  �GD�D$    �D$$�L$��    �L$��L$$��;D�(����   �z43�3�����   ��$    ��u �J03�9,��Ã�;ǋˋ\$|����   �D$�D$�����D$|�����   ���҅��|$ ��   ;|$`�  ���  Uh(�V�� �����7 �D$`PWhd�V� �����\ ��  ����  Uh(�V� ������ �D$�T�@RPh<�V�d ����� �  ����  Uh(�V�A ����� �D$�\�@SSPh��V�! ������ �G  ;|$`u9���9  Uh(�V�� �����n Wh��V�� ����� �  �SP��}(����  Uh(�V� �����. h���~���3���~n�KL�,����q  �D$(;hh�d  �@d��i��   �9h8�D$`��   3ۅ�~���9(��   ����;�|�D$\�\$`9C@��   ��;�|��\$�����[X����A�?  ���M  Uh(�V� ����� �CX���$h��V�� ����� �  ���  �L$\Qh(�V�� �����= UWh\�V� �����f ��  ����  �T$\Rh(�V� ������ UWSh�V�q �����' �  ����  Ph(�V�N ������ �L$`�Q@RUUWh�V�. ������ �T  ���L  �D$\Ph(�V� �����} UWh��V�� ����� �  ��  ���  Uh(�V�� �����< �OH�T$`QRh|�V� �����^ ��   ����   Uh(�V� ������ �GH�L$ PQhH�V�g ����� �   ����   Uh(�V�D ����� �S<Rh�V�+ ������ �T��tPUh(�V� ����� �G(�K<PQh�V�� ����� ��D$`��t�WXRUh��P�� ����q �L$Ld�    Y_^][��D� ��U�l$��L$�  ;iH�  �IDV�D� 9l�(W�<��|$tF�t$ ��t0UhІV�i ������ �W(URh��V�O ����� �@q _^]��� �W43���S��   �O0��    �����*  �D$;XX�  ��k�hxT;_8�|$��   3��~H��9t����;�|��6�D$ 9G@�5  9GD�,  �};�}��9��   ����;�|�|$�D$ 9G@t	9GD�R  ��;���f����|$���_@����A��  �t$$��t4UhІV�^ ������ �G@���$hx�V�@ ������ �1p [_^]��� �|$$��t�UhІW� ����� SVhL�W�� ����� ��o [_^]��� �D$$��t��L$ QhІP�� �L$0���? SWV�t$0Uh�V� hȅV� �� �\����L$$���W���PhІQ� �L$0���� �W@RSSV�t$4Uh��V�^ �D$<�ODPQSh8�V�I ��0�����l$$�������PhІU�) ����� �T$ �GD�O@RPQSSVhȄU� �� ��� ��n [_^]��� �|$$�������UhІW�� �����I �T$�BXPSVh��W� �����j �n [_^]��� [_^�]��� �D$��t�IHQUhP�P�w ���on ]��� ��������U�����E��4S�XxV3���W�xt~l��I ��M���$��|���M�\$8�G���$��|����A�D$8������{8��A��������{R��������At������{���� ;�|��_^[��]������؋E��t�M�Q8Rh�P� ��_^2�[��]����������������������U�l$V3�9w~;�I �G����|&;Ch}!�L$i��   Cd�T$UPQR���������t��;w|�^�]�^2�]���������������V��~ �dot%�F��tj P�po�F    �F    �F    �D$t	V�?������^� ������V��~ �Tmt%�F��tj P�`m�F    �F    �F    �D$t	V��������^� ������S�\$V�3��}^2�[� ��i��   W�yd�8�B@��|k�hAT�xP}_^2�[� �zL U�l$t
�   +U ��U �@L3�90������}	]_^2�[� ��i��   �|8L t�   +�E ]_^�[� ��E ]_^�[� ������������̋T$��i��   V�qd�D0Xk�hAt3ɋp��W~0�x�Ǎ�$    9t
����;�|��|;�}�A�����_^� _���^� ���̋T$��i��   V�qd�D0Xk�hAtW�x�p3�9t�Ǎ�$    ;�}
����9u��|;�}�D1������_^� _���^� ���U����j�h]d�    P��   SUVW�  3�P��$�   d�    �ًCH�sh�L$T�D$<�t$8�d���3����:  �n���3�����    �L$4�Kd݄9�   ��Y`݁�   �Yh�A@��|!݁�   k�hCT���ZX����Au	݁�   �ZX�Sd݄:x  ��:�   �Y`݁�   �Yh�A@��|!݁�   k�hCT���ZX����Au	݁�   �ZX�Cd��X  �D荌8����Y`݁�   �Yh�A@��|%݁�   k�hCT���^X����Au	݁�   �^X�t$8�Kd݄�   ��Y`݁�   �Yh�A@��|!݁�   k�hCT���ZX����Au	݁�   �ZX��   ��������D$4;�}X��i��   +����Kd݄�   �D@ʅ��Y`݁�   �Yh|!݁�   k�hCT���^X����Au	݁�   �^X���   ��u�3�9T$<�T$4�#  �T$8�sDt$8�D$0    �F4���D$@��   �D$0�N0��k�hKT�AX�^@����Au�AX�^@�A<�{$�<�3�9Q@t�   9T�@��   ��Rh�D$DP����U��Ǆ$�       ��v��� ���D$t�$P���*����L$T�P�T$X�H�L$\�P�T$`�H�L$d�P�L$D�T$hǄ$�   �����}� �D$TP�N�`����V@�T$4����Au�^@��؋D$0��;D$@�D$0�����D$8H��;T$<�T$4�������$�   d�    Y_^][��]����������U����j�hS]d�    P��   VW�  3�P��$�   d�    ���wH��蓉����uB���   ��t8�G��|1;��   })i��   ��   ;�u����� ��t;�t
j V���M/ ���F��������D$��   ��\$�F�\$�F�\$$�F�\$,�F �\$4�F(�\$<�} �}�uǄ$�       tU��ti��tM������uBW�L$`�*���PV�L$L����P�L$|�� P�L$Ƅ$�   �C� �L$tƄ$�    ��� ��t�D$��D$�^�D$$�^��t�D$,��D$4�_�D$<�_�L$Ǆ$�   ������ �D$��$�   d�    Y_^��]� ���U����j�h�]d�    P��   SVW�  3�P��$�   d�    �ى\$�L$�� ���   3��Ή�$�   �������   ���   ;�~L�D$���\$���   �|8��8t$�'� �؅�t�L$訇����Q�T$ R���- �Ǩ   �l$u��D$��D$$�^�D$,�^�D$4�^�D$<�^ �D$D�^(���[����؅���   �} ��}�\$�F�\$$�F�\$,�F�\$4�F �\$<�F(�u�\$DtX��tl��tP������uEW�L$P�N��PV�L$l�C��P��$�   ��� P�L$ Ƅ$�   �d� �L$|Ƅ$�    �� ��t�D$��D$$�^�D$,�^��t�D$4��D$<�_�D$D�_�L$Ǆ$�   ������ �Ë�$�   d�    Y_^[��]� �����QS�\$U�l$VW���W83�3��҉T$~(���O4�<� ��t�	��BPSU�Ѕ�tS�T$��;�|ڋW83��҉T$��   ���$    �O$�<� ��t�	��BPSU�Ѕ�tK�T$��;�|�_^][Y� ����   ���$    �O4�<� ��t���BPSU�Ѓ�y�_^]3�[Y� ���t$xL��t$�O$�<� ��t���BPSU��3�9t$~ �O4�<� ��t���BPSU�Ѓ�;t$|��l$y�3�_^][Y� ����������̃�4�T$8S�ً��   V3�;���;�W�D$<�L$�L$�D$ t���:�T$H;�t�2;ƋSx�T$�Sh�T$,�SXU�T$4�t$$�z  �t$���r  ���   D$�x��D$(�9  �H$���L$<}�D$ 3҅ɉT$ �  ��D$(�L$���  �@ ������  ;D$��  k�hCt�H���D$,�L$8}�D$ 3҅ɉT$��  ����$    �D$,�|$ ��  �H�����7  ;T$0�-  �sd��i��   �L0Pƃ����wL�$� J�D$�  �H@����   ;L$4��   k�hKT�yPt
�D$ ��   �yL�;�u�O;�u
�D$ ��   �hLi��   �@X΅���   9D$~�Stk�h�D(���   i��   �|00 t	3�������AX���yL|=9D$~7k�h�L(iɨ   �|10 t	3҅�����t��ta�D$ �Z��uV�D$ �Oh��ḣh7  �1h��ḣh+  � h��ḣhH  �hd�ḣh  hL���b ���T$��;T$8�T$�{����h,�ḣh�  hL��b ���T$ ��;T$<�T$ ������L$�D$$�D$�   ��;D$@�D$$�������u
�D$ �D$ �D$H��]t�T$��D$H��t�T$���t�|$ t�   9��   t���   _^��[��4� �H!H!H@I�T$SV2���W�   ;Qx}zk�hQt�ڋ{��~k3����~c�I ��t\�S����|4;Qh}/i��   Qd�RT��t��t��t��t2���;�|�_^[� h$�h�h�  hL��ea ��2�_^[� ����������3��|$}�Qh�T$W�yh3҅�~+S�\$V3�U;D$}�id9\.<u�������   ;�|�]^[_� �������3��|$}�Qh�T$W�yX3҅�~(S�\$V3�U;D$}�iT9\.<u������h;�|�]^[_� ����������3��|$}
���   �T$W���   3҅�~5S�\$V3�U��$    ;D$}���   9\.,u�����ƨ   ;�|�]^[_� �������QSUV�ًChW�|$�o�O�D$�1 3���~-�O����|;D$}�Sdi��   �����   �҃�;�|�_^][Y� ����������L$�QX����At�|$ u�yP}�QX�	�5�YX�YX����Az�� 2�� �QV��FX����L$~;S�\$UW3���d$ �FT��SP�Bh���Є�u�D$��h��u��D$_][^Y� ��^Y� �������������SV�t$�^(W������ۉN(|F;_H}AU�n4��x7�F0����|(;GX}#k�hGT9X@u�H@9XDu�HDj P����D  �����y�]�F0��t�N8��Qj P�}C
 ���5�F4    _�^@^[� ���̃�S3�U�l$���   �U8;ӉL$�T$�E8������  ;Qh��  �E@;�VW�C  ;AX�:  �t$ k�hAT;��t%�Pu�GL9u�OH������L$VW�6D  �  �EP�wP3҃���3ۃ�����ÉT$�������   ���    �OL��;L$u�WH�B�OHV�ЃP uq���_X�j���}���|`��|\�T$;Jh}S��i��   Bd9H8uC�T$���|�xPu���u�L$�)�D$��������|�xPu�PX;UXu�����t��������T$�d����L$��|�Id3�������i��   �DP���|�Adi��   �DP   3ۋEX;�|6�L$;Ax}-k�hAt���w��x�O�T$9�u�G�P�OV�҃�y�_^�5����U`���   �Uh�E<ݕ�   �E@ݝ�   �ED�EH�EL �]P�]T�EX���   �� S�͉��   �z� ][��� ��QSUV3�W�|$���   9_(�o�l$�G����|	jj�����;���   ;nx��   �_���Fh�D$x6�l$�O����|;D$}i��   FdUP���@X�����d�����yҋl$�G(��|=;��   }5i��   ��   �؋s$��x��    �S 9,�u�C�P�KV�҃�y�3ۉ_$�G;�t�O ��QSP�\@
 ���_�O0�G(������� �_`_^][Y� ������������UV��W���   �ж �|$3퉮�   �G���;ŉO|I;��   }A�FxS�_$���D$x0�l$�W ����|;D$}k�hFtU�H(P�����������y�3�[�O,�G ;�t�O(��QUP�?
 ��U�ωo$��� �OH���   �9� _^]� ���U����j�h�]d�    P��l  SV�  3�P��$x  d�    ��ڋO���L$4��   �G��T$L�P�T$P�P�T$T�P�T$X�P�I�T$\�PɉT$`�ɋT�T$d�T�T$h�T��T$l�T�T$p�T��L$H�T$t�D��L$dQ�L$P�D$|�T����T$|��4������Au��2���$x  d�    Y^[��]���D$4���T$<~G������D$8   �D$D���    �W�؋D$8H�P�����D$<�D$8�l$D�T$<u��D$|���p&������At��L$LQ��$�   R���o���D$dP��$�   Q���o���T$dR�D$PP��$�   �5� �G���S�P�K�H�S�P�K�H�S�L$H�P�G��D��N�H�V�P�N�H�V�P�N�H�D$4�����Ǆ$�      ��   ����   �D$4�G�T$<R�P��$�   ��� �D$<�O��$�   R����$�   �$P�4��n�����d$L��P��$0  Q��$�   R����$(  �$P�n����P��$  Q����m������m�����H�N�P�V�H�N�P�V�@���l$4�F�M�����$�   Ǆ$�  �����R� ���$x  d�    Y^[��]������������U�l$W�}�΋��������U ���   ���ĉ�K�H�K�H�K�H�K�H�K�H���ҋ�U ���   ���ĉ�N�H�N�H�N�H�N�H�N�H����_]���̋T$3���|;QX}k�hQT��� ������V���� ��u���   ��t�v,��|;q8}�A4��^�������V���� ��u;�V`��t4�N<��|-;J(}(�B$�4���th`�hD�h-  hL���V ����^��������V���8� ��u>���   ��t4�N<��|-;J}(�B�4���th��h��h�-  hL��V ����^�����S�\$V��FW�~;�uq��    ��   v��|�  ;�}�������   ~� �V��t.��+���x%;�}!;��}Q���k����V�F���F_^[� ;�}Q���L����N��V_���F^[� �������V��~ ��t%�F��tj P���F    �F    �F    ^�����������VW�|$��;�tB�G��_�F    ��^� 9F}P�tC���N��t�G�F�W�@��PRQ�>
 ��_��^� �����������V��~ ��t%�F��tj P���F    �F    �F    �D$t	V�_�������^� ������j�h�]d�    PQSVW�  3�P�D$d�    �ى\$3�9{8�s,�|$��$t�F;�tWP����$�~�~�~���D$�����	�  �L$d�    Y_^[��������̋A(��}"�L$��tPh��Q�e� ���]R ��� VW�y43���~�Q0�2��|����;�|�_^��  �L$��tVPh`�Q�� ���R _��^� �������������VW3�W���� �5�ԉ����N8�N<�~L�~P�~T�FH�$�^X�~`3��F0�F4_�ND�N@��^�������j�h(^d�    PQSVW�  3�P�D$d�    �ى\$3�9{T�sH�|$��$t�F;�tWP����$�~�~�~���D$�����ɧ �L$d�    Y_^[���������j�hq^d�    PQSUVW�  3�P�D$d�    ��t$耥 3ۃ���~p����n8�n<�n@�^L�^P�^T�nX�\$ �Tm�_�_�_���   �D$ �J� �5ݖ�   3�ݖ�   ���   ���   �F0�F4�Vh�nH�^`�nD�G�   ;��D$ }F9o~�o�O��PUQ����;ÉGt#�O;�}��+���R���SQ��6
 ���o��_�_�ƋL$d�    Y_^][��������������j�h�^d�    PQSVW�  3�P�D$d�    ���|$���   �D$   �� 3�9_|�wp�\$�Tmt�F;�tSP���`m�^�^�^���D$������ �L$d�    Y_^[������j�h�^d�    PQVW�  3�P�D$d�    ��t$�� 3��������F�|$�F�$�~�~�~ �N0�D$�~$�F(譫 3��~`�F�F�ƋL$d�    Y_^�����������������j�h_d�    PQSVW�  3�P�D$d�    ���|$�O0�D$   �� 3�9_ �w�\$��$t�F;�tSP����$�^�^�^���D$�����i �L$d�    Y_^[��������̋Q`��t,�D$��|$;A}�I��3���|;Jh}i��   Jd��� 3�� ��������j�h>_d�    PQSV�  3�P�D$d�    ��t$3�S��� ������F�\$�F�$�^ �^$�^(�NH�D$�F,�^0�^4�I� h@h`�jj�FxP�D$,�r[
 ���   ���   ���   ���   �`/�N8�d/�V<�h/�F@�l/�ND�^�^�ƋL$d�    Y^[�����������j�h�_d�    PQSVW�  3�P�D$d�    ���|$��jj�D$$   蟙��jj��蔙��jj��艙���w3�9^t�F;�t�SP�B���Љ^�^�^h@jj�OxQ�D$,�Z
 �OH�D$�Щ 9^�\$��$t�F;�tSP����$�^�^�^���D$������ �L$d�    Y_^[��������U����j�h�_d�    P��h  SVW�  3�P��$x  d�    ��t$@��P0j�D$H   �ҋ]���]����j �ˉ|$L������\$T��t
ǆ�       ���   �� �^(3���~1��$    �F$�<� ��t� �M��RDQ���҅�u�D$D��;�|֋F8���D$P�D$8    �V  �|$8�F4��ǃ8 �+  3�9\$H��   � ��ȋ��   S�Ѓ�us�N4��P���   �Ѓ�u]�F4�8�Q�� ����tH��� ��V4��؋���   ���$S�҅�u��t��M��PDQ���҅�u��Pj����3ۋF4���E�RDP�҅�u'��t�D$8P�����O������i  �D$D    �\  3�;��R  ��RlW�D$`P���ҋ�Plj�L$pQ�ˉ�$�  ��Ƅ$�  �|$<����   3��d$ W�L$p�X�����D$<P�L$`�X������\$��$�   � �$Q���i �D$8�T$@�r4��W�L$p��^X���D$L�D$<P�L$`�LX���L$L�����\$��$�   � �$R� �D$|P��$�   ��v����;����At�����Q�����L$8Q�L$D���/�����3ۋD$<�����D$<������t��Bj���ЍL$lƄ$�   膦 �L$\Ǆ$�  �����r� �t$@�D$8��;D$P�D$8������FH��~%3��؋ND�9�E�RD�P�҅�u�D$D��H��uߋFX��~3��؋��E�NTP��Һ����h��uꋶ�   ����  �D$T�D$<    ��t$H�\$T�L$@���   \$<�UR��荺���KH�ե ����� ���D$8u$���   ��t\�C,��|U;A8}P�I4�����D$8tB�L$8��$�   R�� ��   �{H󥍌$�   �i� �{�t�L$@�CHP���   蠨 ��4�u�\$T����tXj���3����������DzDj���������X����Dz/j���
������X����Dzj����������X�D$7 ����D{�D$7�|$8��u�D$7 ���   ��tP�|$7 t;W�;�����t1�{0 t9���   �x0��~,3������   �I,���\������u�����   ��BDV�Ѓ��    ��   �|$7 u9��u�    ��$�   �ݔ$�   ݔ$�   ݜ$  ��$�   �`�����tE�L$8Q���   蛞����t1�{0 t<���   �z0��~/3������   �H,��0\������u�����   ��E�RDP�ҋ��   ��tX�|$7 t>�D$8P�:�����t0�{0 t=���   �y0��~03�����   �J,���[������u�����   �M��PDQ���ҁD$<�   �l$H�z����E�L$@P�����D$D��$x  d�    Y_^[��]� �������SV�t$�����W��t[��P4���҃�t5h��h��h  hL��G ��Pt��j���ҋ�P4���҃�u�w�D$P�O����_��^[� _^��[� �������������SV�t$�����W��t[��P4���҃�t5hP�h8�h7  hL��9G ��Pt��j���ҋ�P4���҃�u�w(�D$P�O ����_��^[� _^��[� �������������V��L$W�����t��P4�҃�u�~8�D$P�N0�E������   �
� ��_ǆ�       ^� ���������j�h�_d�    P��SUVW�  3�P�D$$d�    ��l$4�EX3�;���   ;Fx}}�Ntk�h�D(;�|o;��   }gi��   ��   ���������;�tN�E<;�|G;F}B�V�4�;�t8�D$P���� ����   �D$PV�ω\$4�ҍL$�ET��D$,�����$� �ËL$$d�    Y_^][��� ������������QSU�l$�]W�3��ۈD$~DV���    �E�4�i��   qd�|$ t�~P uj V�������FPu�D$��;�|ʊD$^_][Y� ��������������U����j�hm`d�    P��  SVW�  3�P��$�  d�    ��t$$�FX�~�V(�N8�^H�D$8�Fh�D$4�Fx�D$,���   ���|$�T$ �L$0�\$(�D$HuG9D$8��   ����   �E��th�P��� ���B ����$�  d�    Y_^[��]� �|$8 u�E��t�h؟�|$, u�E��t�h��뭅�u�E��t�h��뛃|$4 u�E��t�h��놅�u�E��t�hp��q�����u�E���k���hT��X�����u�E���R���h8��?���3���~H�VD�ʋy(���u)�y4 ~+�U���$����I4QPh�R��� ������;���   ����H;�|�3�9\$8��   �\$�FT�L$�<�G8���u~�P �  9G<�  ����� ���3  ���9G@�F  9GDtS�E��������ODQSh��P�L� �������M���w���P�4��T�(RPh\�Q�$� ���Z���;��  �D$h��;\$8�V����]3�9|$4�J  �|$�Fd�L$ȋA8���;��  9Q@�~  9QX��  9Q<��  9QD��  9QH��   ��������QHRWh�S�� ��������E��������WPRSh��P�p� �������E��������O<QSh`�P�M� �������E���x���Sh�P�.� ���d����E���Y����W@RSh��P�� ���A����E���6����NT��k�h�T
8SRSh��P��� ������;���   ��BS�Ѕ��  �D$�   ��;|$4������T$,3Ʌ��)  �Ft���    �x�����   9x(�v  �x ��   ��������PRQh8�S�Y� ��������������I@QWh��S�9� ���o������g����QXRWh��S�� ���O������G����A<PWh0�S��� ���/������'����IDQWhؚS��� �������������Nd��i��   �T8WRWh��S�� ��������������Wh��S�� �������;���   ����h;������3�9\$H��   �\$�����   �T$�D
����<
��   9G,��  ���� ����  9G$~v9E�^����W$�ERSh8�P�� ���C������;����@(PQh��S��� ���#����������Vt��k�h�DQPQh��S��� �������;��e  �D$�   ��;\$H�>���3�9\$~m�V�<�    �< �tQ� �M��RQ���҅��S  �F���B4�Ѓ��\  �F�8�Q�� ����t���" ���X  ��;\$|�3�9\$ ~m�V$�<�    �< �tQ� �M��RQ���҅��<  �F$���B4�Ѓ��E  �F$�8�Q�� ����t���5" ���A  ��;\$ |�3�9|$0~B�V4�<� ��t-� ��]�ȋBS�Ѕ��,  �N4����B4�Ѓ��2  ��;|$0|�3�9|$(~,3ۋND�|(�t�URW���������   ����H;|$(|�3�9|$8~,3ۋFT�|8�t�MQW���v������  ����h;|$8|�3�9|$H~:3����    ���   �|�t�EPW����������  ���è   ;|$H|�3�9T$,�T$��   �Ft�D$�x�tw�H(���C  ;��   �7  ���   ��i��   9L��  �P3Ʌ҉T$ ~;�P�����  ;Fh��  �^d��i��   9D8��  ����;L$ |̋D$�T$����h;T$,�T$�D$�g���3�9T$4�T$D�T$��	  �T$�~d|$�8���	  �GD����  �NH;���  �GH����  ;��  �GD�ND��9D�(�p
  �GH��9D�(��
  �G<���/  ;F�&  �N�<� ���D$�z
  �GX����  ;Fx��  �Nt�Ћ�k�h9T�x
  �T$k�h�D(�i��   ���   �T$�T,�F4����tS��$�   Q���� �L$����   ��$�   PQ��Ǆ$�      ��9GT�7
  ��$�   Ǆ$�  ������� �P��  �@���  �E��������O@�T$QRhh�P�� ��������} ������G,�MPSh�Q�u� �������E�������Sh��P�V� �������} ��������   ��iɨ   �D�MSPSh��Q�!� ���W����E���L���Sh`�P�� ���8����M���-���PSh,�Q��� �������E������Sh �P��� ��������E�������Sh��P�� ��������M�������PSh��Q�� �������E�������Sh��P�e� �������������Wh`�S�I� �������˅��u���PWh,�Q�*� ���`����E���U���Wh�P�� ���A����E���6���Wh�P��� ���"����E������Wh̖P��� �������} �����QR�Uh��R�� ��������} �����P�D$Q�MPhh�Q�� �������} ������T$P�EQRh8�P�]� �������} �����QR�Uh�R�;� ���q����G@���~	  ;FX�u	  ��k�h^T9C8��  �GL3Ʉ���3҄���OD;L�@����  �WH;T�@��  ��$4  �cL����$L  �WL����$�  �KL����$�  �?L����$d  �3L����$  �'L����$  �L����$|  �L����$�   �L����$�   ��K����Ph��$�   Q����j ��$�   Ǆ$�     �D��� j j ��$l  Q��$@  R�����$����j��$�   �lD��� j j ��$$  Q��$X  R�����$�y����GX�L$$k�hAt�ыp(i��   ��   ���$� ���D$u ���   ��t�v,��|;p8}
�@4���L$݄$<  �t$j j ��$�  R��$  P��$  Q���\$��݄$X  �$�� ݄$T  j j ��$�   R��$�   P��$�  Q���\$��݄$p  �$�R� ��$|  ��Q���Oh��$  �\$<�Q���O`��$�   �D$<�\$L�Q���Oh��$�   �\$<�Q���O`��$|  R���D$H��$�  ݜ$�   ݄$x  �$P��L��݄$t  ��P��$�  Q��$  R����$�   �$P�L��������K����$�  �UQ��݄$$  ��$�   Q����$�   �$R�sL��݄$,  ��P��$�  P��$�   Q����$�  �$R�EL�������kK����$�  ��P����Ph�L$tQ����3�8OLƄ$�  ��Q���9B��� ����$D  �$R�������L$tƄ$�  �� ��Ph��$�   Q����3�8OLƄ$�  ��Q����A��� ����$\  �$R���Q�����$�   Ƅ$�  荐 ��$<  P��$�  �	K���\$<��$T  Q��$�  ��J���D$<�L t��������ɋOD;OHu,�C@;CDu$;�u ����������A�   ��������  ����؍�$  �D$   ��    ���YH�����l$y$�   R��������3�8OL���I���  �P���  �Q�P�Q�P�Q�P�Q�@�A��$�   Q�������3�8OL���I���  �P���  �Q�P�Q�P�Q�P�Q�@�A��$�  Q��$  �;_���\$<��$�  R��$(  �#_���CX���D$L��݄$�   ������'�p&������Au������D$<������A�2  �����������Y  �ٍ�$�   ��Ǆ$�  �������Î ��ܗ�   ����D�V  ܟ�   ����D�v  �]W��~������������Pu�T�G����|  �$����D$D�t$$�T$�D$�   ��;T$4�T$�!����|$, �D$    �d  �D$    �T$$�Zt\$�D$9C�&  ���S@����D�<  �[X����D�\  3�9s�D$ �����D$0�����D$(�����D$������  �K�<��T$$i��   zdj ���   P�K0詎 ���p  j ���   Q�K0萎 ���W  ���U  �S��OD�D$ �L$0�M  �} �o����ERh�P�"� ���X����} �N����MRh��Q�� ���7����} �-����<WWR�Uh��R��� �������E�������ʋT$QRhX�P�� ��������M��t�T$P�GTPRh(�Q�� ���/ ��$�   ��Ǆ$�  ����蟌 �Ƌ�$�  d�    Y_^[��]� �} ������D$�MPh�Q�8� ���n����} �d���V�WL�D$�MRPh��Q�� ���C����} �9���P�����؋E��t%�L t�T$Rhp��
�L$Qh �P��� ����. ��$�   ��Ǆ$�  �����ً �Ƌ�$�  d�    Y_^[��]� �E�م�����t#�T$���\$�\$�$Rh��P�d� ��$�������돋E��t�L$���\$�\$�$Qh`�P�2� ��$�b����E�؅��[���݇�   �T$���$Rh$�P�� ���7����E���,���݇�   �L$���$Qh�P��� ��������� ����T$Rh��S�� ��������E��������O@�T$QRht�P�� ��������} ������MPRhH�Q�i� �������} ������MPRh�Q�G� ���}����} �s����MPRh�Q�%� ���[����} �Q����MPRh��Q�� ���9����T$(;WD��  �C���H��;s�L$�|$(�4����|$  |
9|$0��  �D$�D$h��;D$,�D$������t$$h@h`�jj�T$dR�_:
 3�9D$HǄ$�     �D$0��  �D$ �	��$    ���D$$���   D$ �x �D$,�J  �T$$���O,�B4�4����3  ��Rlj ��$�   P���ҋ�L$T�P�T$X�H�L$\�P��$�   �T$`�#� ��Plj��$�   Q���ҋ�L$d�P�T$h�H�L$l�P��$�   �T$p�� �$ �D$    ~U�G �L$����|1�T$$;Bx}(�Mk�h��CtQ�T$hR�L$\Q������������  �D$�T$,��;B$�D$��|���菐�����D$�I  ����   j ���ҋ�����   j�Ή|$@�҅��D$@u���  �D$�p�L$t�t$�M9����Ƅ$�  �D$    ��  �L$�Q�D$�4��L$$i��   qd�~P�t$L��  �FT���  �|$< �  �x��X��<  �E�؅�������C@�T$���$Rh��P�t� �������E��������CX�L$���$QhL�P�H� ���~����} �t����WD�C���D$R�T$,Q�L$VR�UP���VQhАR�	� ��$�?����E���4����L$VQh��P��� �������} �����T$0�D$ �L$(R�T$P�D$j Q�MR���VPhАQ�� ��$�������u�|$< t�x�X��,��u�|$@ t�x����P  �|$@ �E  �   3�S��$�   R�Ή|$0��������D����$�   S��$�  P���L������eD����$�   ����\$��$�   � �$�DI����t��t�L$t��8����u��   �L$t�_8������   3�;t$��   �T$�B�<��L$$i��   yd�T$(;WTu~�PuxS��$�   P����������C��� ���L$|�$�=7���%�$���5����At;S��$p  Q����������C��� ���L$|�$� 7�����5����A�T  ��;t$�K����D$��;D$�D$�&����L$tƄ$�  �*� �D$0�D$ �   ��;D$H�D$0�}����t$$3�9D$D�D$�E  3ۍ�$    �D$;D$4�.  �Nd���9|8�  �|P��  �D@�l$D��|;D$8|�U���0  k�hFT�D$     �PP�҉T$L��  �PL�T$��I �D$�;T$t.��|*��i��   ��x8�t�xPu�@X;DXu����	  ���D$ �T$L�D$9T$ |����2  ;|$4�(  �DT������F  �$����E��t*�O8�T$LQ�J8�T$ Q�J�T$4Q�JQh��P�� ���& �L$t��Ƅ$�  迃 h@jj�T$`RǄ$�  ������3
 �������i��   �|T��   �E��t�T$WRh��P�A� ���9& h@j��j�D$`PǄ$�  �����3
 �j�����i��   �|
Ttj�E���G  �L$WQh0�P��� ���.  ��i��   �|Tt7�E���  �L$WQhЎP�� ����   ��i��   �|
T��   �D$���   �|$D �����h@jj�D$`PǄ$�  ������2
 �   ��$�  d�    Y_^[��]� �D$Ph��R�9� ���1% ��$�  h@jj�L$`Q���2
 �f����ER�T$WRh@�P��� ����$ Ǆ$�  ����뻋E��t,�L$WQh��P��� ����D$�MPh��Q�� ���$ h@jj�T$`RǄ$�  ��������1
 ������I �x�x�x�xc�����0����̋D$��SUW����   �|$��|y�\$��wpk�hETV��9|�@t�|�@�UD�D$��P�L�,�׫���NP3҅ɉL$~3�FL����|"i��   Ed�xL t	�   +���ˉ|�D�L$��;�|�^_]�[� _]2�[� �����̃�U�l$V3�;�W����  9t$(��  �D$ �t$S��    �D$=   ��  ��~;l$(u����  ��i��   Gd�xPux�L$,�   +މHH�HDU��t�c����輷���   +�;D$(��l$�t$u����   �Odi��   �|P��   �T$R�D$P���h�������   �D$�   �xL �H@t	�   +���ƋT$,RPQ���d�������  ��U��t�ж����)����   +΅����l$�t$��  �Wdi��   xPtP�P@���l  �xL t	�   +���΋wT��k�h�D0P��|StC�L$Q�T$R��譵�����/  �t$�l$�D$��������!�|$ u[_^�]��� �D$,PQR�������D$(�Wd��i��   уzP�D$�D$    uw�D$   ��;D$(t�wd�T$,�T1D�wd�T1HP���0���;D$(t�Wd��i��   �|PtȋOd�D$i��   �t@�����   �L$,3�8PLQ�ϋ�PV������r@����   �GTk�h�|P��   �T$R�D$P��覴�����(  �\$��t�L$Q���:�����T$R��茵������  ��i��   �   +�_dÃxP�l$�t$tf�H@����  �WT��k�h�|*Pu+�xL t	�   +���ƋT$,RPQ���I���[_^�]��� �D$P�L$Q����������~  �l$�t$��l$(�t$ �D$    �^  �d$ �D$=   �K  ��~;l$(u
;t$ �7  ��i��   ÃxPum�L$,�   +މHH�HDU��t�2����苴���   +�;D$(��l$�t$u
;t$ ��   �_di��   �|P��   �T$R�D$P���5����   �xL �H@t	�   +���ƋT$,RPQ���>�������   ��U��t誳��������   +΅����l$�t$|f�_di��   ÃxPtH�P@��|N�xL t	�   +���ƋwT��k�h�L1P��|,t6�T$R�D$P��菲����t�t$�l$�D$�������[_^2�]��� �L$,QPR������[_^�]��� _^2�]��� ����̃��D$P�T$R�D$    �D$   �n�����t�<$ t�|$ u����2�����V���   ��t-��t#��t������t�   ^�ǆ�      3�^Ã��^ø   ^���������������U����j�h�`d�    P���   SVW�  3�P��$�   d�    �L$8��u�V@����At
�} ��  �~4���|$T}�V@�  �5�L$\�^@�\$,�W3���L$<�,���N(3�;���$   �L$(�D$��  ��u�V0�D$������  �L$8k�hAT���ω|$�Ԥ ����  ��Rh��$�   P���ҋ�L$<�P�T$@�H�L$D�P��$�   �T$H�dz 3��_@�D$(9u@V�L$@�}+��� ����$�   �$Q�������MP���J���T$,����Au�\$,��؃�����|��GP3ۅ��D$P�\$$��  �WL�4�����  �D$8;ph��  i��   pd��  ����� ��uK���   ����  �F<����  ;A��  �I�<� ��  h��h��h�-  hL��: �����   ���V  �FX���K  ;Ax�B  �Qtk�h�D(���0  ;��   �$  i��   ��   ���������D$X�  �G@�D$    �   �D$ �d$ �L$(9��   �~L ��u�|$��Rh�D$tP����W��Ƅ$  ��)��� ����$�   �$P���#�����L$\�P�T$`�H�L$d�P�T$h�H�L$l�P�L$t�T$pƄ$    �yx �D$d�L$X���\$��$�   �D$l�$P�v� �MP���:H���T$,�|$����Au�\$,��؋D$ �D$��������D$ �����\$$��;\$P�\$$�����D$��;D$T�D$������;�u�D$,��������Az4�����4�L$<Ǆ$   �����w 2���$�   d�    Y_^[��]� � ��L$<�^@Ǆ$   �����w ���^@����Az����$�   d�    Y_^[��]� ��������������U������l��SV�u�V`W�L$����At�Vh����At
�} ��  �FX����  ;Ax��  k�hAt3ɋx���y  �^8�P9t����;�|��`  �X�D9�����A�4���������?  ���7  �D$�Hh;��(  ;��   �@di��   i��   ���Ћ΋��r����ϋ��i����M�D$�]�������   ����   �|$ ��   �D$P��趾���]�L$0Q���'����T$HR��蛾���D$`P��������3���`�����At�} uvV�؍L$�4��V�L$4���4���� V�L$L���\$��3��V�L$d����3���� ���D$������u�������;������z
� ����������������������l������u�V`����Az�^h����Az�_^[��]� ��_^2�[��]� ̃�SU�l$�E8�ك����V�D$�M8�  ;CX�  W�}P��xk�����EL����|W;Ch}Ri��   Cd���FX���N@|3;Cx}.k�hCt�@(��|!;��   }�L$ i��   ��   QP������j V��跺����y��U@�T$�D$   �I �D$� ��|p;CH}k�SD���t�4���<�x�G0�L$9�u�W,�B�O,V�Ѓ�y�|$  t5�4 /�8 �w,t�F��t�j P�B����3��F�F�FW��薹���D$�l$�v������_�M<�M@�MD�EL3�;�t�MT��QVP�Q�	 ���5�uPV�]X�͉u`�g� ^][��� ��������������j�h�`d�    P��SUVW�  3�P�D$0d�    �ًk8�틳�   �D$�t$$�l$�r  �L$(萵 �EP�L$,�D$<    �;� ����    Q�������j W��	 3���;��D$ ~t�D$���   D$���9Hu�H,�D�@,;�t=��|;�}����u�D$ �����!hD�h(�h"  hL�� ���D$ �D$�   ��u��D$ ��u�K0�����   ;���   3�3�9l$~;�<� t�,����$�S4����t	��Pj�ҋC4��    ��������;t$|ŋt$$3ҋ��   �L,�|;L$}���H,�¨   ��uًt$���x�<� }�S0�B�K0V�Ѓ�y�L$(�D$8������� �S8�K0R�����D$�L$0d�    Y_^][��(����j�had�    P��SUVW�  3�P�D$0d�    �ًk(��sX�D$�t$$�l$�d  �L$(賳 �EP�L$,�D$<    �^� ����    Q�������j W���	 3���;��D$ ~l�D$�CTD$���9H8u�H<�B�@<;�t;|;�}����u�D$ �����!h|�h`�hJ"  hL��� ���D$ �D$h��u��D$ ��u�K �����   ;���   3�3�9l$~;�<� t�,����$�S$����t	��Pj�ҋC$��    ��������;t$|ŋt$$3ҋCT�L<�|;L$}���H<��h��uߋt$���x�<� }�S �B�K V�Ѓ�y�L$(�D$8�����(� �S(�K R�<����D$�L$0d�    Y_^][��(�����j�h8ad�    P��SUVW�  3�P�D$0d�    �ًk��sh�D$�t$$�l$�t  �L$(�� �EP�L$,�D$<    莲 ����    Q�������j W���	 3���;��D$ ~o�D$�CdD$���9H8u�H<�B�@<;�t;|;�}����u�D$ �����!h��h��h�"  hL��� ���D$ �D$�   ��u��D$ ��u�K�߿���   ;���   3�3�9l$~;�<� t�,����$�S����t	��Pj�ҋC��    ��������;t$|ŋt$$3ҍ�$    �Cd�L<�|;L$}���H<���   ��u܋t$���x�I �<� }�S�B�KV�Ѓ�y�L$(�D$8�����H� �S�KR�\����D$�L$0d�    Y_^][��(����̃� S�\$(U�l$0;�V���D$ u'h��hؠhV%  hL�� ��^]2�[�� � �C(��W��  9E(��  �M43����D$�L$,�|$��  ��E0�����D$(�|  k�hFT�H@;M(�D$ u�S(�P@�HD;M(u�S(�PD�PP3Ʌ҉T$$�L$�0  ���D$ �@L���ۉ\$��   ��i��   ~d�OD;M(ut�T$4�B(S�ΉGD腤��3��|X;�tT��   }L��i��   Nd�y@ };�YD�T$8;Z(u
�\$4�[(�YD�YH;Z(u
�T$4�R(�QHP���2����\$����}��l$8�GH;E(uk�L$4�Q(S�ΉWH詣��3���|S�I ;�tL��   }D��i��   Nd�y@ }3�QD;U(u
�T$4�R(�QD�QH;U(u
�T$4�R(�QHP���W�������}��L$��;L$$�L$������\$4�|$�D$(P�K,�Ɩ���L$,��;��|$�c����5�[@����D{
j S�������},3��E(����9_t�G;�t�SP�B���Љ_�_�_U���E����D$_^][�� � �������U����j�hhad�    P��lSW�  3�P�D$xd�    �ً�P4���҃��m  j���]�����A P�L$8�D$,�f 3�9|$(��$�   ~�d$ �L$4����PW���R����;|$(|�U�ˍ|$4������uk�M�9����   ���ĉ8�y�x�y�x�y�x�y�I�x�H���ҋ����   ���ĉ�K�H�K�H�K�H�K�H�K�H�����u���A?��3�9|$(�D$'~b3ۀ|$' ���\$,tW���?���T$,�D$8����$��#���L$8�RW���8P���|$' t�D$,���$W���O������;|$(|��|$@ �D$4�$Ǆ$�   ����t�D$8��tj P�L$<��$�L$xd�    Y_[��]���j�h�ad�    P��,UVW�  3�P�D$<d�    ��l$L���>������u-j ��� ����  VUP�  ���L$<d�    Y_^]��8��T>����P�L$��d �D$$3�P�ˉ|$H�e���P�L$�������$>����~,�L$$QW���s� ��輱��P�L$����˃���=��;�|ԋ΋Ս|$������ul�M ����   ���ĉ�M�H�M�H�M�H�M�H�M�H���ҋ����   ���ĉ�N�H�N�H�N�H�N�H�N�H�����   3��ˉ|$�j=����~v�D$P���� ���td�L$��PRPU�   �D$$���L$$Q�͍t�۰�����H�N�P�V�H�N�P�V�@�F�t$���ˉt$����<��;�|��|$  �D$D�����D$�$t�D$��tj P�L$��$�L$<d�    Y_^]��8��U������4  S�]VWS�XG ������ts�M�9����   ���ĉ8�y�x�y�x�y�x�y�I�x�H���ҋM�9����   ���ĉ8�y�x�y�x�y�x�y�I�x�H����_^[��]�S�} ������  ����   ���҅���   �E�uP����!������  ��$�   Q��������$�   R��$�   P���[!����$�   �o&����4����A�`  ��$@  蒧����$�   Q��$D  讫����RD��$@  P����_^[��]�S谾 ����t�u�]P�]�����_^[��]�S�:������t�MQ�M��������_^[��]�S��� ����t�U�MR���C�����_^[��]ÍD$(P�������L$@Q��葮���uV�L$,�6����4�}����zW�L$D��5����4�����  �D$@P�L$,��5���\$XW���5���T$`����'���D$X����������  ��������A��  �L$@Q��$�   R�L$0�����$P���D$t�$P�r ����W��$�   Q�������$P����$  �$R�E �����D$hP��$,  Q��$  �����$(  �$����4����Au1��$@  �ĥ����$(  R��$D  ������PD��$@  Q���ҍ�$�   P���������L$(�P�T$,�H�L$0�P�T$4�H�L$8�P��$�   P�ˉT$@������L$@�P�T$D�H�L$H�P�T$L�H�L$P�PV�L$,�T$X�U4����4��������Au!��W�L$D�84����4��������A�M  �D$`�d$X��������A��   �D$@P��$�   Q�L$0�6����$P����$  �$R������L$x�P�T$|�H��$�   �P��$�   �H��$�   �P����$@  �T$|�k����D$`�t$X�L$h�T$l�� ���\$���$�   �P��$�   �H��$�   �P��$�   �H��$`  �P�������PD��$@  Q���ҍ�$�   P���)�����L$(�P�T$,�H�L$0�P�T$4�H�L$8�P��$�   P�ˉT$@�q�����L$@�P�T$D�H�L$H�P�T$L�H�L$P�PV�L$,�T$X�2����4��������Au!��W�L$D�2����4��������A��  �\$`����A��  �D$hP��$�   Q��$  �����$P����$�   �$R�Z������$�   P��$�   Q�L$0�����$�   ��!����$�   R��$�   P���{����$�   ��!����$�   Q��$�   R��$�   P��#������$�   �c!���T$X��4������   ��$�   �!����$�   P��$�   �>���\$`��$�  �^����D$`��$�   ��$�   ���ĉ��$�   �P��$�   �H��$�   �P��$�   �H��$�   �P��$�   ���ĉ��$�   �P��$�   �H��$�   �P��$�   �H���P�\$݄$�   ��$   �$�ݪ����PD��$�  Q����������؋����   ���ĉ�N�H�N�H�N�H�N�H�N�H���ҋ����   ���ĉ�O�H�O�H�O�H�O�H�O�H����_^[��]�������̃�|U�o`����  S��������؅ۉ\$��  V�D$@P���.����D$H�L$@�T$D�D$0�D$T�D$<�G@���L$(�L$L�T$,�T$P�L$4�T$8|N�UD���ʍ4ʋPj ���҅�t5�D$pP���G����L$(�P�T$,�H�L$0�P�T$4�H�L$8�P�T$<�D$XP�������D$`�L$X�T$\�D$�D$l�D$$�GD���L$�L$d�T$�T$h�L$�T$ |N�UD���ʍ4ʋPj ���҅�t5�D$pP���G����L$�P�T$�H�L$�P�T$�H�L$ �P�T$$�D$@P�L$,�������^t�G@��|�UD�5���\�@2ۍD$TP�L$�����t�GD��|�UD�5���\�@���u �T$�5�D$�_XP�L$(QR������[]��|������j�h�ad�    P��DSUVW�  3�P�D$Xd�    ��|$h���D$ ��  ;}X��  k�h}T�z  �8 �p  �����������_  ��Ph�L$8Q���ҍD$(P���D$d    �Z ��Rh�D$P���D$d�ҋ��D$`�Y ����   �D$(P�L$<�?%������   �D$p����   }�O<jQ���{�������   �T$8R�L$�%������   �G<�M$�T$���	���ĉ�T$,�P�T$0�P�T$4�P�l�����tX�L$�T$���ĉ�L$0�P�T$4�H�ωP��X �L$�T$���ĉ�L$0�P�T$4�H�ωP�Z\ �D$��   ���i1������t ����   �L$(Q���҅�u?��Pj���ҍL$�D$`��\ �L$(�D$` ��\ �L$8�D$`�����\ 2���   ���HX ��t����   ���҅�t��L$�T$���ĉ�L$0�P�T$4�H�ΉP�m�����Ph�L$HQ���ҍL$Q���D$d�#���L$H���D$`�>\ ��t��Bj�����G���V���r���V�ωG<�y �L$�D$`�	\ �L$(�D$` ��[ �L$8�D$`������[ �|$ t�|$l t�g����D$�L$Xd�    Y_^][��P� �������������j�h bd�    P��@SUVW�  3�P�D$Td�    ��|$d2ۅ��l  ;}h�c  i��   }d�T  �8 �J  ���@��������9  ��Ph�L$4Q���ҍD$$P���D$`    ��W ��Rh�D$P���D$`�ҋ��D$\�V ����   �D$$P�L$8�O"������   �O<jQ���J�������   �T$4R�L$�#"������  �G<�M�T$���	���ĉ�T$(�P�T$,�P�T$0�P苏����tS�L$�T$���ĉ�L$,�P�T$0�H�ωP�V �L$�T$���ĉ�L$,�P�T$0�H�ωP�yY ��   ���.������t ����   �L$$Q���҅�u?��Pj���ҍL$�D$\��Y �L$$�D$\ ��Y �L$4�D$\������Y 2���   ���lU ��t����   ���҅�t��L$�T$���ĉ�L$,�P�T$0�H�ΉP葎����Ph�L$DQ���ҍL$Q���D$`�� ���L$D���D$\�bY ��t��Bj�����G���V������V�ωG<��v ��L$�\$\�,Y �L$$�D$\ �Y �L$4�D$\�����Y �ËL$Td�    Y_^][��L� �����U������DSVW���͍���sp3�9~t�F;�t�WP�B���Љ~�~�~���   ;�u2�_^[��]� �S8R�������t��������;���   �M��PDQ���҅�tƍD$ P���� �����   �   �L$ �PX �u��j ݓ�   ��ݛ�   �6����@j �Kh���\$�#���� j�K`���D$�\$�����@j�Kh���\$������{T �C`��D$�D$���[`���[ht���   S�CT    ����_^�[��]� ���������������V��F�V;�u=�@�Ɂ�   v��|���� ;�}�������   ��;�}P���&����N�I�N��3���A�A�N�F�I���N��^�������������j�hQbd�    PQVW�  3�P�D$d�    �t$ �t$3�;��|$t5���n  �5����F(�����F,�$�~0�~4�~8�^@3��F �F$�L$d�    Y_^��� ��j�h{bd�    PQVW�  3�P�D$d�    jH覟�������t$3�;��|$tI����m  �5����F(�����F,�$�~0�~4�~8�^@3��F �F$�ƋL$d�    Y_^���3��L$d�    Y_^���������j�h�bd�    PQSVW�  3�P�D$d�    ��jH���������t$3�;�\$t7���Ym  �5����F(�����F,�$�^0�^4�^8�^@3��F �F$�3�;��D$����t3;�t/W����m  �G �F �O$�F,�@�N$�W(�N,�V(�W,R���G@�^@�ƋL$d�    Y_^[������V�������D$t	V�K�������^� ��j�h�bd�    PQ�  3�P�D$d�    jh�������D$���D$    t��讥���L$d�    Y���3��L$d�    Y���������������j�hcd�    PQVW�  3�P�D$d�    ��jh褝�����D$���D$    t���:������3����D$����tW���<���ƋL$d�    Y_^���������������V���H����D$t	V�;�������^� ��j�h;cd�    PQ�  3�P�D$d�    h�   �������D$���D$    t���k����L$d�    Y���3��L$d�    Y������������j�hkcd�    PQVW�  3�P�D$d�    ��h�   葜�����D$���D$    t����������3����D$����tW���M=���ƋL$d�    Y_^������������V���إ���D$t	V�+�������^� ��j�h�cd�    P��SUVW�  3�P�D$$d�    ��~p3�9_t�G;�t�SP�B���Љ_�_�_��蛇��3�9��   ��   ��Rh�D$P���ҋF8���   P�\$0�������tS���a�����;�tF����   ���ЍL$���D���L$�T$���ĉ�L$,�P�T$0�H�ωP�-���W���o �L$�D$,�����R ;�u����^ ��;�t09^@�FD�NH�FH�ND��|8^L�VL�L$$d�    Y_^][��ËŋL$$d�    Y_^][����������������j�h�cd�    PQ�  3�P�D$d�    jh訚�����D$���D$    t��辤���L$d�    Y���3��L$d�    Y���������������j�h�cd�    PQVW�  3�P�D$d�    ��jh�4������D$���D$    t���J������3����D$����tW���`=���ƋL$d�    Y_^���������������V��蘤���D$t	V�˛������^� ��j�h+dd�    PQ�  3�P�D$d�    h�   蕙�����D$���D$    t�������L$d�    Y���3��L$d�    Y������������j�h[dd�    PQVW�  3�P�D$d�    ��h�   �!������D$���D$    t��藤�����3����D$����tW���=���ƋL$d�    Y_^������������V���8����D$t	V軚������^� �̃�S�\$�CUVW�����   3��9C�t$}P���e���;�~|�l$���   �L$ƃ�t.��t!��t���   ��u$���   ��u���   ����   ����   ��t��4  �D$ �L$ P�������|$  u�D$�ƨ   �l$u�9l$u�C+�x;C�C_^]3�[��� _^��][��� ��������QS�\$U�kV�3���W���D$~0��    �C��i��   Gd��P虬����u�D$��;�|ڊD$_^][Y� ��������������QS�\$U�k$V�3���W���D$~2��    �C ���L$k�hGtQP��������u�D$��;�|؊D$_^][Y� ������������U����j�h�dd�    P��h  SVW�  3�P��$x  d�    �ى\$`�}h��W�z� ���   ����u/��~+���   �x$u�@ � P���O�����thĥW�@� ���C8Ph��W�.� �C(Ph��W�� �CPh��W�� �CHPh��W�� �CXPht�W�� �ChPhd�W�� �Cx��HPhT�W�є ���   PhD�W返 �C�����D$D    ��  ���$    �K�T$D�4����[  ��Ph�L$lQ���ҍL$|Ǆ$�      ������$�   ������$�   P���q�����L$|�P��$�   �H��$�   �P��$�   �H��$�   �P��$�   P�Ή�$�   誔�����$�   �P��$�   �H��$�   �P��$�   �H��$�   �P���$�   ����ҋ��P_������u�k4j�L$p�
���j �L$p�D$L�����݄$�   �L$H�T$D��0�\$(݄$�   �\$ ݄$�   �\$݄$�   �\$��\$� �$VRh�W�L� ��@�L$lǄ$�  �����eK ��D$DPh��W�#� ���D$D��;C�D$D�l����{( �D$D    �q  �K$�T$D�4����8  ��Ph�L$lQ���ҍL$|Ǆ$�     �V����$�   �J����$�   P���˒��� �\$|��$�   �@Qݜ$�   ���@ݜ$�   �"���� �ݜ$�   ���@ݜ$�   �@�ݜ$�   �Ћ���]������u�k4j�L$p����j �L$p�D$L����݄$�   �L$H��@�\$8��$�   ݄$�   �\$0݄$�   �\$(݄$�   �\$ ݄$�   �\$݄$�   �\$��\$� �$VRh��W�ɑ ��P�L$lǄ$�  ������I ��D$DPh��W蠑 ���D$D��;C(�D$D������{8 �D$D    ��  ��$    �K4�T$D�4����a  ��Plj ��$   Q���ҋ�Plj�L$pQ��Ǆ$�     �ҋ���Ƅ$�  �ҋ��\�����D$Tu�D$Tk4j�L$p�^���j �L$p�D$L�O���j��$   �D$`�=���j ��$   �D$h�+����L$H��T$\�L$d�� �\$��T$t�\$��\$� �D$d�$RPh��W萐 ��0�{8u`���   ��uU��~Q���   �x$uE�@ �Q���_�����t4���ԏ h��W�I� ����迏 ��BW���Ћ��� ���� �L$lƄ$�  �FH ��$�   Ǆ$�  �����/H ��L$DQhl�W�� ���D$D��;C8�D$D�f����CH���D$P    ��   �D$L    �sDt$L�T$P�F@�� �\$�F�\$�F�\$�F�$RhD�W膏 ��,�~4 ~x����� h<�W�k� ���~4 �D$D    ~@���$    ��|$D �x:u�t:�N0�T$D��QPW�-� �D$P����;F4�D$D|ʋ��ӎ hKW�� ���D$P�D$LH��;CH�D$P�1����CX���D$P    ��  �D$L    ��sTt$L���FX�V<�FD�$�N@R�T$\PQRh�W褎 �� ���� ����p ��uH�N`���.  �F<���#  ;A(�  �I$�<� �  h`�hD�h-  hL��:� ����$�   R���X�����$  P���Ɏ����Rh�D$lP���҉D$H��Ph��$�   Q��Ǆ$�     �҉D$\�L$HjƄ$�  �D����L$\j �D$L�5���݄$  �L$H��@�\$8݄$T  �\$0݄$L  �\$(݄$�   �\$ ݄$�   �\$݄$�   �\$��\$� �$hԣW�v� ��H��$�   Ƅ$�  �E �L$l�   ��Rh��$�   P���҉D$H��Ph�L$|Q��Ǆ$�     �҉D$\�L$HjƄ$�  �q����L$\j �D$L�b����L$H����\$� �$h��W�� ���L$|Ƅ$�  �E ��$�   Ǆ$�  ������D �FP����   Ph��W裌 ���~P �D$D    ~c���VL�D$D�������|!;Ch}�Sd��i��   �|L ���u��#�|$D ���u���PQRW�B� �D$T����;FP�D$D|�hKW�$� �����ڋ �D$P�D$Lh��;CX�D$P�1���3�9��   �D$L��  �D$P����$    �ً��   t$P�Ήt$H�)n ���D$hu ���   ��t�F,��|;A8}
�I4���T$h�F0�N,�T$LPQRh`�W舋 ���~$ �D$X    ~=��$    �|$X �x:u�t:�N �T$X��QPW�M� �D$d����;F$�D$X|�hKW�/� ����襊 ���   ��th�D$DXf��������D$Tt4h A���J�����u
�D$DPf��L$Th�A�.�����u�D$DHf���   �' �T$DPRh@�W越 �����   ��t�' Ph$�W蘊 ���D$L��|7;��   }/���   D$P�x$u�@ � P���h�����th�W�Y� ���~$ �D$X    �  �d$ �L$H�Q �D$X���L$`��k�hYt�C$���\$\w#�$�(��������آ��̢��,1�KQPRh��W�� 3���9s~'���x:u�t:�S��QPW軉 ����;s|�hKW襉 ������ �{ �D$T    �>  ���$    �T$\�B�L$T�4��T$`��$�   i��   rd���k ���D$du@���   ��t6�F<��|/;A}*�I�����D$dth��h��h�-  hL��� ����$�   ������$�   �����FP��wC�$�<��D$D���:�D$D���0�D$D���&�D$D|���D$Dp���D$D̢��D$D,1�FT��w8�$�T��k4�/�h��(�X��!�H���@���0��� �����Fh�VH�FD�N@���\$�F`�$R��$�   PQRhԡW�0� ��(��覇 �F<�NL�T$DPQSRh��W�� ���|$d ���   ��$�   P�������$�   �P��$�   �H��$�   �P��$�   �H��$�   �P��$�   P�Ή�$�   �E������$�   �P��$�   �H��$�   �P��$�   �H��$�   �P��$�   ��Ph�L$|Q���ҋ؋�Ph��$�   Q��Ǆ$�     �ҋ�j��Ƅ$�  	����j �΋�����݄$�   ��0�\$(݄$  �\$ ݄$  �\$݄$�   �\$��\$� �$h��W�ۆ ��8��$�   Ƅ$�  ��> �L$|Ǆ$�  ������> �|$h �;  ݄$�   �t$h���\$��$  ݄$�   ���$P�ʪ ݄$�   ���\$��$�   ݄$�   �$Q��裪 ݄$�   ��0�\$(݄$�   �\$ ݄$�   �\$݄$L  �\$݄$D  �\$݄$<  �$hX�W�� ��8�   ��Rh��$$  P�ҋ؋�Ph��$4  Q��Ǆ$�  
   �ҋ�j��Ƅ$�  ����j �΋���������\$� �$h4�W蘅 ����$4  Ƅ$�  
�= ��$$  Ǆ$�  �����= ���#� �D$T�L$\��;A�D$T��������� �D$X�T$H��;B$�D$X��������� �D$L�L$`�D$P�   ��;��   �D$L�"�����$x  d�    Y_^[��]� ��������(�2�<�F�P�Z�{�������������V��~` u2�^� SU�n0W����< 3�9~~E�F�����N`|0;Ah}+i��   Ad��t�L$Q��������t�À   S����? ��;~|�_][�^� _][2�^� ������SV��^��xCW�<�����N�9�P�j �ҋFjH�j P�|�	 �Nσ�Q�����������H��}�_�F    ^[��������S�\$��UVW��}N3�9nt:�~��x!����ۋN��P�U�҃���H;�}�N��PUQ���҉n_�n�n^][� �F;�}x�N��PSQ����3�;ǉFtT�V��+ʍ����Q�ҍ�WP��	 �F��;�}"�<������+�N�Q��������H��u�_�^^][� �~�~_^][� ~V���;�|'�<���+������N�9�B�j �Ѓ�H��u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� �����j�h1ed�    P��SUVW�  3�P�D$ d�    ��}���|$��   k�h3ۋ��M�9�P�S�ҋEjh�SP��	 �u����t$�t$�\$(tCS����1 �5����ԉ�N8�N<�FH�$�^L�^P�^T�^X3��^`�F0�F4�ND�N@�����D$����h;ÉL$(�D$�n����]�L$ d�    Y_^][����E    �L$ d�    Y_^][���������������j�haed�    P��SVW�  3�P�D$d�    ���_��xe��i��   ���    �O�1�P�j �ҋGh�   �j P��	 �O��ΉL$�L$�D$     t����������   ���D$ ����}��G    �L$d�    Y_^[����j�h�ed�    P��SVW�  3�P�D$d�    ���_��xT��k�h�O�1�P�j �ҋGjh�j P���	 �O��ΉL$�L$�D$     t�΋������h���D$ ����}��G    �L$d�    Y_^[�����j�h�ed�    P��SVW�  3�P�D$d�    ���_��xe��i��   ���    �O�1�P�j �ҋGh�   �j P�O�	 �O��ΉL$�L$�D$     t而������   ���D$ ����}��G    �L$d�    Y_^[����SW�|$����~dU�l$��|ZV�t$��|P;�tL�C�/;�B;�>�K�>;�~�;�}��P���f����C�����R�L� ��R����R��	 ��^]_[� �����������S�\$��U��~[W�|$��|QV�t$��|G;�tC�E�;�9;�5�M�;�~�;�}��P�������Ek�hk�hk�hS��WV��	 ��^_][� ����S�\$��U��~dW�|$��|ZV�t$��|P;�tL�E�;�B;�>�M�;�~�;�}��P���v����Ei��   i��   i��   S��WV�%�	 ��^_][� �����������S�\$��U��~[W�|$��|QV�t$��|G;�tC�E�;�9;�5�M�;�~�;�}��P���6 ���Ek�hk�hk�hS��WV访	 ��^_][� ����S�\$��U��~dW�|$��|ZV�t$��|P;�tL�E�;�B;�>�M�;�~�;�}��P���� ���Eiۨ   i��   i��   S��WV�5�	 ��^_][� �����������U����j�h�ed�    P��UVW�  3�P�D$(d�    ��3�9n`��   ��Ph�L$Q���ҋF8�N`UUP�l$<�G�����tS���|�������tF����   ���ҍL$�������L$�T$���ĉ�L$,�P�T$0�H�ωP�i��W��� R �L$�D$0�����4 ��u���DA ���th�F@�ND�FD�F`���N@tU�VP���xhxJ�5�FL����|3;�}/�N`i��   Ad�xL ���HL�Hx��~�@t������� ��u��y��؋ŋL$(d�    Y_^]��]��QS�\$U�k$V�3���W���D$~-��    �C ��k�hGt��P������u�D$��;�|݊D$_^][Y� �UW��3�9o�hmt>V�w��x#S����ۋO��P�U�҃���H;�}�[�O��PUQ���҉o^�o�o_]���������QW�����   ����L$~<S�\$UV3��萋��   �SP��������u�D$�ƨ   ��u܊D$^][_Y� ��_Y� ��������̋D$��S�U�V�t$�PV���c���������t)��t%;�t!W3�9{~����B���Ѓ���H;{|��_^][� �����������V��V2���tQ�N��~JW�|$��t@��~9WjHQR��, 3���9~~%S3����    �F���B�Ѓ���H;~|�[�_^� ���������������V��V2���tQ�N��~JW�|$��t@��~9WjHQR�u, 3���9~~%S3����    �F���B�Ѓ���H;~|�[�_^� ���������������UW��3�9o�|mt:V�w��xS��k�h�O��P�U�҃���h;�}�[�O��PUQ���҉o^�o�o_]������������̋D$k�hSUV�t$PV���ɔ��������t)��t%;�t!W3�9{~����B���Ѓ���h;{|��_^][� �V��V2���tQ�N��~JW�|$��t@��~9WjhQR�U+ 3���9~~%S3����    �F���B�Ѓ���h;~|�[�_^� ���������������UW��3�9o��mt:V�w��xS��k�h�O��P�U�҃���h;�}�[�O��PUQ���҉o^�o�o_]�������������V��V2���tQ�N��~JW�|$��t@��~9WjhQR�* 3���9~~%S3����    �F���B�Ѓ���h;~|�[�_^� ���������������V�������D$t	V�z������^� ��V����������D$t	V�z������^� ������������V�������D$t	V�kz������^� ��V��� ������D$t	V�Ez������^� ������������V�������D$t	V�z������^� ��SUV��W�N@�����NP�*������   �����N`�'����Np������^3�3�;�~$�d$ �F��;�t	��Bj�ЋN�,���;�|��F;�t�V��RUP�ڷ	 ���n�N;�t�F;�~��PUQ躷	 ���^(3�;�~ �N$��;�t	��Bj�ЋN$�,���;�|��F$;�t�V,��RUP�x�	 ���n(�N$;�t�F,;�~��PUQ�X�	 ���^83�;�~ �N4��;�t	��Bj�ЋN4�,���;�|��F4;�t�V<��RUP��	 ���n8�N4;�t�F<;�~��PUQ���	 �����   �- _���   ^][�������������̃�0SVW��3��q����|$@�;�t[����D$,�D$0�D$4�D$8�D$�D$ �D$$�D$(�D$P�T$ R�D$4PQ�Ή\$�\$ �\$$�\$(��� ��t�_^�[��0� _^��[��0� �V�񃾤    u2�^� SW3�9~$~6�\$��F �������   |;Ax}k�hAttS���������t��;~$|�_[�^� _[2�^� ���������������VW�|$����|y;~}t�NS����ۋ�P�j �ҋFjH�j P觵	 �N+σ���Q�WRW�������F�NjH���T��j R�x�	 �F�N���T����R��������F�[_^� �����̋D$9A}	�D$������ �����������UW��3�9ot@V�w��x%S����ۋ��O��P�U�҃���H;�}�[�O��PUQ���҉o^�o�o_]�������������V��F�V;�uN��k�h��   v��|�C� ;�}�������   ��;�}=P�������N��k�hF���N^�k�hFj ��ȋB�ЋNk�hNQ���#����N��k�hF���N^�S�\$��V��|u;^}p�NW��k�h�9�P�j �ҋFjh�j P��	 �N+˃���Q�SRS���s����F�Nk�hjh�T�j R�ܳ	 �F�Nk�h�T���R�������F�_^[� ����������S�\$��V����   ;^��   �NW��i��   �9�P�j �ҋFh�   �j P�m�	 �N+˃���Q�SRS���E����F�Ni��   h�   ��8���j R�5�	 �F�Ni��   ��8�����R���7����F�_^[� �������������V��V2���tT�N��~MW�|$��tC��~<Wh�   QR�$ 3���9~~%S3���I �F���B�Ѓ����   ;~|�[�_^� ������������S�\$��V��|u;^}p�NW��k�h�9�P�j �ҋFjh�j P�[�	 �N+˃���Q�SRS�������F�Nk�hjh�T�j R�,�	 �F�Nk�h�T���R�������F�_^[� ����������UW��3�9ot@V�w��x%S��k�h��    �O��P�U�҃���h;�}�[�O��PUQ���҉o^�o�o_]�������������S�\$��V����   ;^��   �NW��i��   �9�P�j �ҋFh�   �j P�]�	 �N+˃���Q�SRS���%����F�Ni��   h�   ��X���j R�%�	 �F�Ni��   ��X�����R��������F�_^[� ������������̋D$i��   SUV�t$PV������������t,��t(;�t$W3�9{~����B���Ѓ��ƨ   ;{|��_^][� �����������V��V2���tT�N��~MW�|$��tC��~<Wh�   QR�! 3���9~~%S3���I �F���B�Ѓ��è   ;~|�[�_^� ������������V��V2���tT�N��~MW�|$��tC��~<Wh�   QR�"! 3���9~~%S3���I �F���B�Ѓ��è   ;~|�[�_^� ������������������������ ����������j ��m�3�������4����������j ��m�������j�h�fd�    PQSVW�  3�P�D$d�    ��t$�1� 3�W�N�|$ ��������W�N �D$ ����W�N0�D$ �� �~D�~H�~L�F@H��~T�~X�~\�FP\��~d�~h�~l�F`p��~t�~x�~|�Fp�����   ���   ���   ǆ�   �����   ���D$�$ �L;��D$	t�3��F�F�ˉ��   �% �ƋL$d�    Y_^[�����������j�hgd�    PQV�  3�P�D$d�    ��t$���jj�D$	   ��0�����   �D$�$ ���   j �D$��m�	����Np�D$�4�������N`j �D$��m�q����NP�D$� ������N@�D$�������N0�D$订 �N �D$葔���N�D$ 脔�����D$�����ŉ �L$d�    Y^�������SUV��W�}H�w9uL�]@}V���������|;s�s�MD�5�����x(����P����H����P����H���_^�P����X@]�H[����������{����D$�L$�X@�T$�H�L$�P�T$�H�L$�P�T$�H�P�  �������SVW���_X�OP�����5���D$�^X���^8�F<|;G(}�O$��R���@ �~`_��^[� ���������j�h@gd�    P�� SUVW�  3�P�D$4d�    ���_X�OP�<����5���D$L�^X�n8�] 3�;ÉF<|;G(}�O$��R���@ �D$D�~`�H(�|$H�N@�W(U�H,�VD��L��U�O,��L���|$P;���   ��������t{�L$�R����D$$P�Ή\$@�� WP�L$�D$D������L$$�\$<�" �L$�L�����t'�L$�T$���ĉ�L$,�P�T$0�H�ΉP� �L$�D$<������! �D$T���^X�L$4d�    Y_^][��,� �SUV��nxW�}�^pǆ�       9{}W���������|;{�{�L$��k�hFt_�p`^�h]�H$[� ��SUV��W�{x�w�kpǃ�       9u}V���z�����|;u�u�D$��k�hst���n�} �|$�F$�^`�O�N(uM�G$����|L;Gu���ab��9G}P���Ժ���G�G���Pj j���>����W�E _��^`��^][� U�O�1K��_�^`��^][� ����̃�0SUV��W���   �  ���   �}���   ǆ�       9{}W���������|;{�{�D$D��iۨ   ��   ���k�C,���   |F;F8}A�N4��R���9 ���>J ��t(�D$P���.J ���7� ���{H�   �L$�� _^]��[��0� ������SW�����   ���~)UV3��苇�   �P��������u2ہƨ   ��u�^]_��[���UV�t$k�hW��wt3�F���D$~;S�I �N���Od��i��   �|
D }���a����P(RS���U����D$��;�|�[_^]� ���j�h�gd�    P��   SUVW�  3�P��$�   d�    ��$�   ��wO���    tF�Wl������t;��PlU�L$(Q���ҍL$$Ǆ$�       ������u2�L$$Ǆ$�   ����� 3���$�   d�    Y_^][�ļ   � ��P0j���ҋF,���   jP�|b����~"��Bd���Ћ��   ��W� |��W�ΉF,��7 ����   U���Ѕ��v����L$$�T$(�D$,�L$�L$0�T$�D$�L$ �L$Ƅ$�   �������RlU�D$8P����P�L$Ƅ$�   �>����L$4��Ƅ$�   �� ��t[�L$�T$���ĉ�L$,�P�T$0�HU�ωP�/o ��PlU�L$8Q���ҋ�L$�P�T$�H�L$�P�L$4�T$ �l j�L$H�A^��j �L$����j�L$���y�������\$�L$D� �$�B�������̉�P�Q�P�@�Q�T$8�A�L$4���ĉ�L$L�P�T$P�HU�L$hƄ$�   �P��t���L$4Ƅ$�   �� �D$DP�������3�9~$~,��N �������   |;Ax}k�hAttP�a����;~$|Հ~0 ���   �V0���   ��t��u
ǁ�       ���   ��tU�������   U�������   ��tU��������   U�����L$Ƅ$�    �" �L$$Ǆ$�   ����� �   �`�������j�h�gd�    P���   VW�  3�P��$�   d�    �񃾤    ��   ��E ����u$���   ��t�F,��|;A8}�I4�<�����   ��B0j���ЋN,jQ���   �_����~"��Bd���Ћ��   ��W�/y��W�ΉF,��4 ��Rlj �D$ P���ҋ�Plj�L$Q��Ǆ$�       �ҋ���   ��Ƅ$�   �҅�u>�L$��$�   � �L$Ǆ$�   ������ 3���$�   d�    Y_^���   Ë�Plj �L$@Q���ҋ�Plj�L$0Q��Ƅ$�   ��j�L$PƄ$�   �x[��j �L$P�\����j ��L$P�~\����j�X�L$P�n\����j��L$P�_\�����X�΍D$LP�^���3�9~$~2��$    �N �������   |;Ax}k�hAttP�^����;~$|Հ~0 ���   �ɈV0t�������   �A������   ��t�������   �'����L$,Ƅ$�   �� �L$<Ƅ$�   � �L$Ƅ$�    � �L$Ǆ$�   ����� �   ��$�   d�    Y_^���   ����j�h<hd�    P��T  SUVW�  3�P��$h  d�    �ك��    Ǆ$p     ��$x  u+Ƅ$p   � ��$�  Ǆ$p  ����� 2��  �F�������  ��$�  �2�������  ���Cf�������  �E �Plj �L$Q���ҋE �Plj�L$(Q��Ƅ$x  �ҍ�$x  P�L$Ƅ$t  �F�����t��$�  Q�L$(�1�������  j��$l  �;Y��j�L$l�0Y��j��$�   �"Y����$x  R�L$������tb��$x  ��$|  ���ĉ��$�  �P��$�  �H�L$$�P�T$(���ĉ�L$<�P�T$@�Hj ��$�   �P�o������  ��$�  P�L$(������tb��$�  ��$�  ���ĉ��$�  �P��$�  �H�L$4�P�T$8���ĉ�L$L�P�T$P�Hj��$  �P�<o�����6  ��$�   P��$�  Q�L$p�[Y������B0�    ��$h  �j���ЋK,jQ���   �[����~#�U �Bd���Ћ��   ��U��t��U�ˉC,�0 �L$Q��$|  �6�����t9��$x  ��$|  ���ĉ��$�  �H��$�  �P�Hj ���-h ��t{�T$$R��$�  ���������   ��$�  ��$�  ���ĉ��$�  �P��$�  �Hj�͉P��g ��uW�L$�T$���ĉ�L$,�P�T$0�Hj �͉P�g �L$$Ƅ$p  � �L$Ƅ$p  �� ��$x  ������E �Plj �L$8Q���ҋ��$x  �P��$|  �H��$�  �P�L$4��$�  � �E �Plj�L$8Q���ҋ��$�  �P��$�  �H��$�  �P�L$4��$�  �n j��$�   �@V��j�L$l�5V����$x  P�L$������tb��$x  ��$|  ���ĉ��$�  �P��$�  �H�L$$�P�T$(���ĉ�L$<�P�T$@�Hj ��$  �P��l�����������$�  P�L$(�-�����tb��$�  ��$�  ���ĉ��$�  �P��$�  �H�L$4�P�T$8���ĉ�L$L�P�T$P�Hj��$�   �P�Ol�����I����D$hP��$�  Q��$�   �nV����    ��$h  ��$h  �R���?������	������   ���   ���   �D$T�L$X�T$\3ۋl�T���Q  3��w������D$$u�D$��P�L$4�H�T$8�P�L$<�T$@����$�  u��$x  ��P�L$D�H�T$H�P�L$L�T$P��Ƅ$p  ���������   �D$DP�L$8���������   �L$4Q���$�����t�T$D��D$H�F�L$L�N�T$P�V�kj ���j���� ���L$<�$�������L$L�$�j����\$`j���=���� ���L$<�$�������L$L�$�=������\$���D$p�$������L$DƄ$p  �� �L$4Ƅ$p  � �������������������L$$Ƅ$p  � �L$Ƅ$p  �| ��$x  Ƅ$p   �h ��$�  Ǆ$p  �����Q ���$h  d�    Y_^][��`  �  ���j�hphd�    P�� UVW�  3�P�D$0d�    ���l$@���+  �5���D$D��������D�  �D$L��������D��   ��������   ���    ��   �_��������   ��Plj �L$$Q���ҋ�Plj�L$Q���D$@    ���D$L�����\$�D$T�D$H�$�L$ u�L$0�d����L$�T$���ĉ�L$(�P�T$,�H�L$0�P�T$4���ĉ�L$H�P�T$L�H�ωP�����L$���D$8 �� �L$ �D$8������ �ƋL$0d�    Y_^]��,� ����3��L$0d�    Y_^]��,� ���������j�h�hd�    P��SUVW�  3�P�D$0d�    ���|$���   3�;��D$�t$ ��  �L$(�R �FP�L$,�\$<�0S ���    Q�E ������SU蕙	 �Wx��3�;�T$$~m�\$�D$���   t$�F���u�D� �8;�u�^�\� ���(hd�hH�h�!  hL�蜴 �N���D$ �L� �D$�   ��;|$ |���u_�l$�ŀ   9]tE�u��x$��i��   �M�9�B�j �Ѓ���   ��}�U �E�Rj P�����E    3ۉ]�]�   �t$ ;���   ���x>��i��   �L$���   �|��DuV���   �������L� �����   ��}ʋ|$$��~L3��T$�Bt�L0(ƃ��|;L$ }	�L� �H(�!h,�hH�h�!  hL�膳 ���D$ ��h��u��L$(�D$8�����R �|$���   ���   R�����D$�L$0d�    Y_^][��(��������j�h�hd�    P�� SUVW�  3�P�D$4d�    ��t$�^x3�;��D$�\$ �  �L$,�DP �CP�L$0�|$@��P ��    Q� ������WP�D$(�W�	 ���   �Fh��3�;߉T$$�D$(~z3�����$    �t$�vt�D���u	�L$���>;�u�T$�n�,����+h�hЧh�"  hL��I� �F�L$,���D$ ������h;|$ |���u�t$�Np�����.  �t$ ;��  ���x7��k�h�l$�Ut�|��DuV�Mp������	�L$�������h��}���l$�D$$��~|3ۉD$$���   �D$�x���|V�F ������|#;D$ }�T$����|��/�F�P�NW���!h��hЧh�"  hL��`� ���D$ ��y��è   �l$$u��|$(��~R3��D$�@d�L0Xƃ��|;L$ }�T$���HX�!h��hЧh #  hL���� ���D$ ���   ��u��t$�L$,�D$<�����P �Vx�NpR�[����D$�L$4d�    Y_^][��,����j�h�hd�    P�� SUVW�  3�P�D$4d�    ��t$�^h3�;��D$�\$ ��  �L$,��M �CP�L$0�|$@�sN ��    Q� ������WP�D$(�ה	 �Vx�FX��3�;߉T$$�D$(~t3���t$�vd�D8���u	�L$���>;�u�T$�n8�,����+ht�hX�h"#  hL��կ �F8�L$,���D$ �������   ;|$ |���ud�t$�~d �n`tJ�u��x'��i��   �I �M�9�B�j �Ѓ����   ��}�U �E�Rj P���ҋt$�E    3��E�E�\  �t$ ;��L  ���x@��i��   �I �l$�Ed�|8��D8uV�M`�����	�L$��������   ��}���l$�D$$���v   3ۉD$$�ut�D�x���|V�F������|#;D$ }�T$����|��/�F�P�NW���!h4�hX�h=#  hL�茮 ���D$ ��y���h�l$$u��\$(���u   3�D$�pT�D.P��x���|W�NL�������|#;D$ }�T$����|��/�FH�P�NHW���!h�hX�hS#  hL��	� ���D$ ��y���h��u��t$�L$,�D$<�����M �Fh�N`P�#����D$�L$4d�    Y_^][��,������������j�h(id�    P�� SUVW�  3�P�D$4d�    ��t$�^X3�;��D$�\$ ��  �L$,��J �CP�L$0�|$@�sK ��    Q� ������WP�D$(�ב	 �VH�Fh��3�;߉T$(�D$$~q3���t$�vT�D8���u	�L$���>;�u�T$�n8�,����+h �h�h|#  hL��լ �F8�L$,���D$ ������h;|$ |���u�t$�NP�G����"  �t$ ;��  ���x7��k�h�l$�UT�|8��D8uV�MP������	�L$�������h��}���l$�|$$��~N3��Ed�L0@ƃ��|;L$ }�T$���H@�!h��h�h�#  hL��� ���D$ ���   ��u��\$(��~t3�T$�rD�D.4��x���|V�F0������|#;D$ }�T$����|��/�F,�P�N,W���!h��h�h�#  hL�虫 ���D$ ��y���H��u��t$�L$,�D$<�����J �FX�NPP�����D$�L$4d�    Y_^][��,������������j�hXid�    P��$SUVW�  3�P�D$8d�    ���|$�wH3�;��D$�t$��  �L$0�TH �FP�L$4�\$D�I ��    Q� ������SP�D$,�g�	 �Gh�WX��;ÉD$,�T$(��   �D$$����    �|$�od�}8���   �}D��|B;�}>�D$�HD�4�����|1(�u'h �h�h�#  hL��R� �T$(�BD���|0(�}H��|D;|$}>�L$�QD�4�����|2(�u'h��h�h�#  hL��� �D$(�HD���|1(�t$���   �l$$�D���3�3���~o3ۋT$�rD�D(���u�D$ �������>;�u�L$ �n(�,����+hl�h�h�#  hL�菩 �V(�D$0���D$ ������H;|$|���u�L$��@������  �t$;��  ���x=�<�������l$�MD�|9(��D9(uV�M@������	�T$ �������H��}���l$�D$(��~^3ۉD$$�ETÍp@�   ����|;D$}�T$ ����!hH�h�h$  hL�辨 ���D$ ����u���h�l$$u��\$,��~_3�L$�AdōpD�   ����|;D$}�T$ ����!h$�h�h#$  hL��X� ���D$ ����u����   ��u��L$0�D$@�����\G �|$�WH�O@R�l����D$�L$8d�    Y_^][��0�����j�h�id�    P��(SUVW�  3�P�D$<d�    �ى\$�D$�Y���3��u�D$��������u�D$���i�����u�D$���j�����u�D$���������u�D$���������u�D$���͐����u�D$��莒����u�D$�D$�H�l$ �l$$�l$(�s�Kh;�l$D�*  ��~V�L$ �BC���l$ ���D$(|;��t$$��t��~Pj U蝋	 �l$,��3҅��~F3�����   �Kd�9Q8u�I<��|;�}�<) u
�)�l$ �2������   ;�|Ą���   3�;��D$,�D�D$0�D$4�D$8~V�L$0��-���l$ 3Ʌ�~.3ҋCd�k�|<�|� �l$0|� �H<�����   ;�|؋l$ 3Ʌ�~�T$0���C����;�|�l$ �|$8 �D$,�Dt�D$0��tj P�L$4��D�l$ �s(;sX��  �D$(;�~y��~R9t$$~�t$$�D$�PVU�L$$�ҋ�3�;�l$ t#�L$(;�~��+�RP�Q�S�	 �l$,���t$(�-�D$(�D$$�#��t�D$�P3�WU�L$$��3�l$ �|$(�|$$��|
;t$(�t$$��t�|$( ~�D$(Pj U��	 �l$,��3҅��~E3�������   �KT�9Q8u�I<��|;�}�<) u
�)�l$ �2�����h;�|Ǆ���   3�;��D$,�D�D$0�D$4�D$8~V�L$0�+,���l$ 3Ʌ�~+3ҋCT�k$�|<�|� �l$0|� �H<����h;�|ۋl$ 3Ʌ�~�D$0���S$����;�|�l$ �|$8 �D$,�Dt�D$0��tj P�L$4��D�l$ �s8;��   �   �D$(;�~y��~R9t$$~�t$$�T$�BVU�L$$�Ћ�3�;�l$ t#�L$(;�~��+�RP�Q誈	 �l$,���t$(�-�D$(�D$$�#��t�D$�P3�WU�L$$��3�l$ �|$(�|$$��|
;t$(�t$$��t�|$( ~�D$(Pj U�J�	 �l$,��3҅��~I3����@  ���   �9Qu�I,��|;�}�<) u
�)�l$ �2����Ǩ   ;�|����  3�;��D$,do�|$0�|$4�|$8~V��}�t$4Vj �L$4�po�����|$0t)�D$8;�~��+���Q��j R蝇	 �|$<���t$8�
3��D$8�D$4�l$ 3҅�~<3����$    ����   �[4�l,��ȉ��\$�Q,�|$0���   ;�|ԋl$ 3Ʌ�~���C4���|$0��;�|�l$ �|$8 �D$,dot"��t3�VW�L$4�po�l$ �t$0�t$8�t$4�|$( �D$D�����D$�Ht��tj U�L$$��H�D$�L$<d�    Y_^][��4��j�h�id�    P��4SUVW�  3�P�D$Hd�    ��\$X;���  �&���S���b �CH�u@P�������CX�}PP����������   ���   P�`����Ch�M`P������Cx�MpP�����CH��|;F�F�CX��|;G�G���   ��|;��   ���   �Ch��|;El�Eh�Cx��|;E|�Ex�EP�K�s���M Q�K �s���U0R�K0�P{ �MH��~Y3��D$X�L$�sD�}D��;�t3V���y  �F �G �N$�G,�@�O$�V(�O,�W(�V,R���F@�D$X�_@��H�l$�D$Xu��EX���B  3��D$�{T�MT��;��L$XtFW�� �O0�D$X�H0�W4�P4�O8�H8�W<�P<�O@�H@�WD�HH�PD��@�WHR���GX�L$X�YX�}T�D7<����o`|�U$���D$X��D$X    �KT�T$�R��� ����̉�P�Q�P�@�Q�A�L$hQ���D$d    �u �L$�D$P������ �KT��� ��t���� �ST��@h��T$(R�Ћ���̉�P�Q�P�@�Q�A���D$`   �� �L$(�D$P������ ��h�l$������Mx��~3��Ut�l`��h��u񋅈   ���r   3��t$X�D$���t$X���   ���   �P��������   �D7,������   |�M4���3�P���� ���   �D$X�   ��H�l$�tH�   �u��Eh���   3��D$�Cd�Md�P�������}d�D7<������   |�M���T$X��D$X    �Kd�D$(�P�T� ����̉�P�Q�P�@�Q�A�L$hQ���D$d   �� �L$(�D$P�����t� �Kd��
� ��t���/ �Sd�2�@h�2�T$8R�Ћ���̉�P�Q�P�@�Q�A���D$`   �b� �L$8�D$P������ ���   �l$�����Mx���l   3��D$X�L$�st�}t��;�tFV������N�O�V�W�F�W�R�O�G�FP�ҋF$�G$�N(�D$X�O(��0��0�   ��h�l$�D$Xu����   ���   �   󥋓�   ���   �ŋL$Hd�    Y_^][��@� ��V��F�V;�u@��i��   ��   v��|�x=
 ;�}�������   ��;�}2P�������(i��   Fj ��ȋB�ЋNi��   NQ���[����N��i��   F���N^������V��j ��m������D$t	V��B������^� ����������V���4������D$t	V�B������^� ������������V��j ��m������D$t	V�cB������^� ����������j�h�id�    PQ�  3�P�D$d�    h�   �%@�����D$���D$    t��������L$d�    Y���3��L$d�    Y������������j�h+jd�    PQVW�  3�P�D$d�    ��h�   �?�����D$���D$    t���w������3����D$����tW�������ƋL$d�    Y_^������������VW�|$��t5h�P���:����t%�t$��th�P���"����tW������_�^�_2�^�������������j�h[jd�    PQ�  3�P�D$d�    h�   ��>�����D$���D$    t�������L$d�    Y���3��L$d�    Y������������V�������D$t	V�@������^� ��j�h�jd�    PQSUVW�  3�P�D$d�    ��t$�l$(U�Z 3�W�N�|$$����Ve��W�N �D$$�He��W�N0�D$$�Js �~D�~H�~L�F@H��~T�~X�~\�FP\��~d�~h�~l�F`p��~t�~x�~|�Fp�����   ���   ���   ǆ�   �����   ���D$ ��� �L;��D$ 	t�3��F�F�ˉ��   �w� U�������ƋL$d�    Y_^][��� ������̃�0SUV��W�~h3ۍN`���   ������5��D$D�U`����Uh;�ݕ�   ݝ�   ���   �}8�M@�]P�]L�E<�]T�MX���   |I;F}D�N�4�;�t:V���W �T$R����] �����   �   �L$�� ��ݕ�   ݝ�   _^��][��0� ��������̋D$VWPǁ�       �*����|$�O8���V8�N@R�OH�����D$3Ʌ����T�@3Ʌ������VD���T�@�FL_�VH��^� ���j�hkd�    P��4SUVW�  3�P�D$Hd�    �ًD$X�t$d�T$\Vǃ�       �HPR�L$P���P����l$`���E�O8Q�M�|$h�GX�D����|t;s}o�S�4���te�L$��� j �D$P���D$X    �B] ��t1�}���T$(�\$@u�}0�   �t$�|$d��L$Q�M0�� �L$�D$P�����<� �t$��u	�GP   �y��u'�T$X�BL�i��   Kd�AX+E������GP�AP�M3҅��D$d   ~8�L$X�[d�m�IL�d$ �i��   �9hXt����;�|���   �HP�L$d�T$d�WP�ǋL$Hd�    Y_^][��@� ����������j�hHkd�    P��0SUVW�  3�P�D$Dd�    ��|$\Wǆ�       �����|$T �l$X�����CL�M�S8�KXR�M������|p;~}k�F�<���ta�L$�t� j �L$Q���D$T    �[ ��t-�}���T$$�\$<u�}0�   �t$���T$R�M0�� �L$�D$L������ �ËL$Dd�    Y_^][��<� ���̋D$�T$PRj �������L$�I(�P`�T$�Phݐ�   �HDݘ�   �HH�@P   �PTǀ�   	   � ���U����j�h{kd�    P���   SUVW�  3�P��$�   d�    ��l$X�UX���   �����~3���I �ET���h���p@�pDu�Uh��~3ɍd$ �Ed����   ���pD�pHu�u@���p����FP���ų���EX+��   ���� }�    9F}P��袳����~E�D$8    �|$<�����   |$83��_$��~�O ��R���������;�|�D$8�   �l$<uɋuH�L$d�t$D虧���L$|萧��3�;��|$8��  �|$<�L$d������}D�\$\|$<3ۋG4���D$@�P  ��$    �G0������   k�hET���~< ��   ���� ��uH�N`����   �F<����   ;A(��   �I$�<� ��   h`�hD�h-  hL��@� ���D$89F@u��$�   R���U6���9FDuS��$�   P���6��� �T$|�@ݔ$�   �@ݔ$�   �D$d�����\$d�D$l�\$l�D$t�\$t�D$\��$�\$\��;\$@�������D$\��������AuD��L$d��Q����$�   �$R�Ѩ����O�P�W�H�O�P�W�H�O�P���W��؋D$8�D$<H��;D$D�D$8�o���3��uX�ƙ�������3�;ǉt$D�D$H��|$L�L$P�|$T~P�L$L�����L$P;���$   ��   3ۋuT�D@����   �ND��|;�t{���J ��u8�N`��ti�F<��|b;A(}]�I$�<� tTh`�hD�h-  hL�衑 ������   ���Ѕ�t(�L$H�����ND�V@;�}
��ND�H���V@�P�x����h;|$D�Y����L$P����  �D$L��t#�`��t��~h`jQP��� �L$`�������|$D�D$@   ��   ���    ���D$7 ��   �T$L�   �D$<3�|$8;ǋ*�\*}=�u+�92�2u��T$L�D$79Xu��P��T$L�D$7����uЋ|$D�D$<�����l$8�D$<u��|$7 �L$Pt>��t'��~#�`��t��~h`jQR�(� �L$`���D$@��;ǉD$@�>���3����D$7 ��   �t$L�@�ҋ<2�X;�}�,[�4��d$ ;>u
����;�|�;Ë�}V��+ȋ�L$@���L$L�D);�~0����|*;�}&�T$X;rH}�ʋAD����R����P��|���D$7���l$@u��L$P;ً��m����|$7 t	�L$X�L����|$T Ǆ$   �����D$H�t�D$L��tj P�L$P����$�   d�    Y_^][��]�������j�h�kd�    PVW�  3�P�D$d�    ���t$��t;�tHW��������3h�   �\3�����D$���D$    tW����������3��D$����jj�������ƋL$d�    Y_^��� ��V�t$��th�Q���������t��^�3�^���������������̸�Q�����������S���׫���؄�u�D$��th��P�^1 ����[� ����V�t$WhܫV���=1 ����W���4 h�&V�$1 ��_^� ������������VW�|$j ��j����4 ����t��V���1 ��_^� ��̃�VW�|$��D$P�L$Q���D$    �D$    ��4 ����t�|$u��V��� ��_^��� VW�|$W���r���W��Vjjj j��� ��_��^� ����̋D$�T$PR��Qjj蹻 ����� j�h�kd�    PQV�  3�P�D$d�    ��t$�M ����T$�T$�N�$�D$,    ���=����ƋL$d�    Y^�������������V���XM �D$����N�P�V�H�N�P�V�H�N�P�V��^� ��������uM �����VW�|$��;�t-W�>M �O�G�N�P�V�H�N�P�V�H�N�P�V_��^� j�hld�    PQ�  3�P�D$d�    j �h0�����D$���D$    t�������L$d�    Y���3��L$d�    Y���������������j�h;ld�    PQVW�  3�P�D$d�    ��j ��/�����D$���D$    t���J������3����D$����t3;�t/W���<L �O�G�N�P�V�H�N�P�V�H�N�P�V�ƋL$d�    Y_^����VW�|$��t5h�Q���Z�����t%�t$��th�Q���B�����tW���v���_�^�_2�^�������������V������K �D$t	V�1������^� ������������V�t$��tI���f= w*f=0 r7f=9 vf=A r+f=Z vf=_ tf=a rf=z wf��0�Srf��9w���2�^�2��V����f�� rf��"tf��tf��0r�f��9r���f�> u��uf�~� w2�[^���������j�hhld�    PQV�  3�P�D$d�    ��t$���  ���   �D$    �����ƋL$d�    Y^����������������j�h�ld�    PQV�  3�P�D$d�    ��t$���   �D$    �������D$�����&�  �L$d�    Y^��������V����  �D$t	V�/������^� ��VW�|$W����I �G�F�O�N�W�V�G�F�O�W�NR�N��/ �G �F �O$�N$�W(�V(�G,�F,�O0�N0�W8�V8�G<�F<�O@�N@�WD�VD�GH�FH�OL�NL�WP�VP�GT�FT�OX�NX�W\�V\�G`�F`�Od�Nd�Wh�Vh�Gl�Fl�Op�Np�Wt�Vt�Gx�Fx�O|�N|���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ݇�   ݞ�   ݇�   ݞ�   ݇�   ݞ�   ݇�   ݞ�   ݇�   ݞ�   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ݇�   _ݞ�   ��^� ���������������V��N� �F    諑��ǆ�       ��^��������������SV�񋆸   3�;�t 9v� ����   9wP�y-�������   9��   u�N;�t8t	��Pj�҈�^^[�������������j�h�ld�    PQV�  3�P�D$d�    ��t$�D$    �k����N�D$�����;����L$d�    Y^�������������VW�|$W������G�F�O�N�W�V�G�F�O�W�NR�N�H- �F �P�N �� W��_��^� ��SU�l$V2���� ��9��  t.��t�D$Ph��U�) h�U�	) �����  ^]�[�^]��[����̋D$� �L$+���̋L$��T$+u�A+B������������j�h�ld�    PQSUVW�  3�P�D$d�    �ى\$�l$(U�1 �EP�K�D$$    ��0 �u�{�	   �u,�{,�	   �MP�KP�ËL$d�    Y_^][��� ��������������̋T$��@j Rj j ��3Ʌ������ ��S�\$UVW��   �Wh(�S�D. �u ���˃��& P����Ѕ�|������ |�h �����, _^][� �����������S�\$UVW��   �Wh<�S��- �u ���˃� �$& P����Ѕ�|������ |�h4����, _^][� �����������VW�|$��;~tjS3�;�~I9~~�~�N��PWQ����;ÉFt?�V;�~��+ʍ���Q����SP�h	 ��[�~_^� �F;�t�SP�B�Љ^�^�^[_^� ���̋Q2���t%�I��~V�t$��t��~VjQR�x� ���^� ��������������̋Q2���t%�I��~V�t$��t��~VjQR�(� ���^� ��������������̋D$�T$��    QR�
B����� ���̋Q2���t(�I��~!V�t$��t��~Vh�  QR��� ���^� �����������̋Q2���t(�I��~!V�t$��t��~Vh�  QR�� ���^� �����������̋Q2���t(�I��~!V�t$��t��~Vh�   QR�U� ���^� �����������̋Q2���t(�I��~!V�t$��t��~Vh�   QR�� ���^� �����������̋D$�L$�@��PQ��@����� ����̋Q2���t%�I��~V�t$��t��~Vj0QR�� ���^� ��������������̋Q2���t%�I��~V�t$��t��~Vj0QR�h� ���^� ���������������VW�|$W�������GP�N�f( �O�G�N��V�H�N�P�V�@�F_��^� ���������������SU�l$VWU���@����EP�K�( �M�K�U�S�E�C�E�[�M �K �U$�S$�E(�C(�M,�K,�U0�͉S0�C4+˺A   ��f�4f�0����u񍵸   ���   �   󥋅  _^��  ]��[� ���������VW�|$W�������GP�N�v' �O�N�W�V�G�F�O�N�W�V�G �^ �G(�^(�G0�^0�G8�^8�G@�^@�GH�^H�GP�FP�OT�NT�WX�VX�G\�F\�O`�N`�Wd�Vd�Gh�Fh�Ol�Nl�Gp�^p�Wx�Vx݇�   ݞ�   ���   ���   ���   ���   ���   ���   ���   ���   Q���   ���   �& ���   R���   �& ���   P���   �& ���   Q���   �s& ���   ���   ݇�   ݞ�   ݇�   ݞ�   ���   ���   ���   ���   ���   _���   ��^� ���j�h1md�    PQ�  3�P�D$d�    �L$�L$���D$    t�&� �L$d�    Y��� ����j�hamd�    PQ�  3�P�D$d�    �L$�L$���D$    t�F�  �L$d�    Y��� ����j�h�md�    PQ�  3�P�D$d�    �L$�L$���D$    t�v� �L$d�    Y��� ���̋Q2���t(�I��~!V�t$��t��~Vh�  QR��� ���^� �����������̋Q2���t(�I��~!V�t$��t��~Vh�  QR�� ���^� �����������̋D$�L$i��  PQ�{<����� �����j�h�md�    PQ�  3�P�D$d�    �L$�L$���D$    t���  �L$d�    Y��� ���̋Q2���t(�I��~!V�t$��t��~Vh�   QR��� ���^� �����������̋Q2���t(�I��~!V�t$��t��~Vh�   QR�� ���^� �����������̋D$�L$i��   PQ�;����� ����̋D$�L$�@��PQ�k;����� �����j�h�md�    PQ�  3�P�D$d�    �L$�L$���D$    t�j �L$d�    Y��� ���̋Q2���t%�I��~V�t$��t��~VjpQR��� ���^� ��������������̋Q2���t%�I��~V�t$��t��~VjpQR�� ���^� ��������������̋D$�L$k�pPQ�~:����� �������̋Q2���t%�I��~V�t$��t��~Vj QR�H� ���^� ��������������̋D$�L$��PQ�:����� ��������j�h!nd�    PQ�  3�P�D$d�    �L$�L$���D$    t�� �L$d�    Y��� ���̋Q2���t(�I��~!V�t$��t��~Vh  QR�� ���^� �����������̋Q2���t(�I��~!V�t$��t��~Vh  QR�E� ���^� �����������̋D$�L$i�  PQ�+9����� �����j�hQnd�    PQ�  3�P�D$d�    �L$�L$���D$    t�vG �L$d�    Y��� ���̋Q2���t(�I��~!V�t$��t��~Vh�   QR�� ���^� �����������̋Q2���t(�I��~!V�t$��t��~Vh�   QR�U� ���^� ������������j�h�nd�    PQ�  3�P�D$d�    �L$�L$���D$    t�&U �L$d�    Y��� ���̋Q2���t%�I��~V�t$��t��~Vj8QR��� ���^� ��������������̋Q2���t%�I��~V�t$��t��~Vj8QR�� ���^� ���������������j�h�nd�    PQ�  3�P�D$d�    �L$�L$���D$    t�&� �L$d�    Y��� ����j�h�nd�    PQ�  3�P�D$d�    �L$�L$���D$    t�v	���L$d�    Y��� ����j�hod�    PQV�  3�P�D$d�    �t$�t$���D$    t7�`/��d/�N�h/�V�l/�N�F�Q� �F(    �F,    �L$d�    Y^��� SU�l$VWU�������E�C�M�K�U�S�E�C�M�U�KR�K�F �E �C �M!�K!�U$�S$�E(�C(�M,�K,�U0�S0�E4�C4�M8�K8�U<�S<�E@�C@�uH�{H�    󥋍�   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ݅�   ݛ�   ݅�   ݛ�   ݅   ݛ   ݅  ݛ  ݅  ݛ  ��  ��  ݅   ݛ   ݅(  ݛ(  _݅0  ^ݛ0  ݅8  ݛ8  ��@  ��@  ��D  ��D  ��H  ��H  ��L  ��L  ��P  ��P  ��T  ]��T  ��[� ���������̋D$� V����H�N�P�V�H�N�P�V�H�N�P�V�H �N �P$�N(��(�V$�P�B�Ћ�^� ̃��|$ W��tF3��D$�D$�F���L$t1�N��~*h &jQP�D$P�&t	 ����t�N+�����|�|���|;|$|	�D$_��Ë�_�����̋A8�QVP�AR���   �L$P�s�����^� �����������̋A<�Q VP�A	R���   �L$P�C�����^� ������������V��~ ���t%�F��tj P����F    �F    �F    ^����������̋D$�L$����PQ�3����� ����SW�|$����~bU�l$��|XV�t$��|N;�tJ�C�/;�@;�<�K�>;�~�;�}��P�������C����R�L� ��R����R��X	 ��^]_[� ������������̋A@�Q$VP�A
R���   �L$P�3�����^� ������������V��L$��|9�F;�}2+���P�APQ���,����F��N�V3�������A�A�A�A^� ��������QSW�|$j �ً�PWj j �\$�҅�}��th��W� ��_2�[Y� V�t$����   ��|H�� ;�?��2|�gfff������������+�u�P��� �ȸgfff���������;�~43���t.��� P�� �ȸgfff���������QVhP�W�| ��U�l$����� ��u ���h
  h�W�V ��]^_2�[Y� �K�1���PV���O ��u ���3
  h�W�! ��]^_2�[Y� �SR���	� ��u ���
  h��W�� ��]^_2�[Y� ���   S���w� ��u ����	  h�W�� ��]^_2�[Y� ���\� �؄�u ����	  hȸW� ��]^_2�[Y� 3��d$ �D$;��  }4���  ����Q��� � �؄�u��tVh��W�J ������u������ ��u ���4	  h@�W�" ��]^_2�[Y� ���	  ���� ����   ���F� �؄�u"�ǅ���  h��P�� ��]^_2�[Y� 3�3����$    ��T$;��  }?���  �P���"� �؄�u�|$$ t�L$$Wh��Q� �����Ƹ  ��u����μ ��u$�D$$���e  h`�P�S ��]^_2�[Y� ���E  ���Ǽ �؄�u$�D$$���,  h�P� ��]^_2�[Y� 3�3����$    �T$;��  }?���  �P���� �؄�u�|$$ t�L$$WhжQ�� �����Ƙ   ��u����N� ��u$�D$$����  h��P� ��]^_2�[Y� ����  ����� ����   ���w� �؄�u$�D$$���\  hL�P�J ��]^_2�[Y� 3�3����$    �T$;��  }<���  �P���"� �؄�u�|$$ t�L$$Wh �Q�� ������0��u����� ��u$�D$$����  h��P�� ��]^_2�[Y� ����  ���z� �؄�u$�D$$����  h��P� ��]^_2�[Y� 3�3��T$;��  }<���  �P���� �؄�u�|$$ t�L$$Wh@�Q�A ������p��u����m� ��u$�D$$���$  h �P� ��]^_2�[Y� ���  ��膹 �؄�u$�D$$����  hĴP�� ��]^_2�[Y� 3�3����    �T$;�   }<���  �P���b� �؄�u�|$$ t�L$$Wh��Q� ������ ��u����� ��u$�D$$���h  h@�P�V ��]^_2�[Y� ���H  ���� ����   ���ڸ �؄�u$�D$$���  h�P� ��]^_2�[Y� 3�3��T$;�  }?��  �P���N� �؄�u�|$$ t�L$$Wh��Q�� ������  ��u����j� ��u$�D$$����  h��P� ��]^_2�[Y� ����  ����� ����   ���3� �؄�u$�D$$���X  hD�P�F ��]^_2�[Y� 3�3���I �T$;�   }?��  �P���2� �؄�u�|$$ t�L$$Wh��Q�� �������   ��u���辷 ��u$�D$$����  h��P�� ��]^_2�[Y� ����  ���׻ �؄�u$�D$$����  h|�P� ��]^_2�[Y� 3�3����$    �T$;�0  }G��,  �1���   RP����� �؄�u�|$$ t�D$$Wh8�P�- �����Ɛ  ��u����V� ��u$�D$$���  h��P�� ��]^_2�[Y� ����  ���_� ����   ��迶 �؄�u$�D$$����  h��P� ��]^_2�[Y� 3�3���L$;�@  }<�ы�<  �P���B� �؄�u�|$$ t�D$$Wh`�P�e ������8��u����Q� ��u$�D$$���H  h�P�6 ��]^_2�[Y� ���(  ���� ����   ���:� �؄�u$�D$$����  hȰP�� ��]^_2�[Y� 3�3��L$;�P  }?�ы�L  �P���� �؄�u�|$$ t�D$$Whx�P� �������   ��u����ʵ ��u$�D$$����  h0�P�o ��]^_2�[Y� ���a  ��裹 �؄�u$�D$$���H  h�P�6 ��]^_2�[Y� 3�3���I �D$;�`  }T��\  �|1 t:�Ћ�\  �T0ƍHQR����� �؄�u�|$$ t�D$$Wh��P�� �������   ��u����� ��u$�D$$����   hl�P� ��]^_2�[Y� ����   ���� ����   ���� �؄�u �D$$��tkh(�P�Y ��]^_2�[Y� �|$3���    ;�p  }��l  ����t
P���S� �؃���uڋ�蓴 ��u �D$$��th�P��
 ��]^_2�[Y� ��t���D$    tT3����$    �d$ �T$�D$;��  }5�ʋ�|  �V��#������t�F,�N(�VRPQV���� �D$��0뻋��$� ��u�D$$2ۅ�th��P�k
 ��]^_��[Y� �������������̃�,�  3ĉD$(�D$0�T$8SU�ًL$<V�L$(�D$$�D$H�L$$WQ�T$4�D$8�D$�����:#��������  ��`  ���t$��  ���  ��谳 ;��a  ���1� V���Y� 3����H  3����$    �d$ ��\  �L�D�L$�P�T$�H�L$ �P�D$P�T$(�"������tKh<�h$�h�  hH��Of �L$(Q������\  �L$,�D��T$0�P�L$4�H�T$8���P�L$�T$jW���ĉ�L$8�P�T$<�H�͉P�� ��uuh�h$�h�  hH���e �D$(P�|����\  �T$,�D��L$0�H�T$4���P�L$$j �H�T$�L$ W���ĉ�T$8�H�L$<�P�H���� �����   ;|$������L$(�T$R�T$0���ĉ�L$D�P�T$H�H�͉P�K� ��u���_^][�L$(3��E	 ��,� �L$8�D$_^][3��E	 ��,� �����̃�,�  3ĉD$(�D$0�T$8SU�ًL$<V�L$(�D$$�D$H�L$$WQ�T$4�D$8�D$������ ��������  ��P  ���t$��  ���  ���p� ;��a  ���� V���� 3����H  3����$    �d$ ��L  �L�D�L$�P�T$�H�L$ �P�D$P�T$(�? ������tKh��hp�h�  hH��d �L$(Q�����L  �L$,�D��T$0�P�L$4�H�T$8���P�L$�T$jW���ĉ�L$8�P�T$<�H�͉P��� ��uuhT�hp�h�  hH��c �D$(P�<����L  �T$,�D��L$0�H�T$4���P�L$$j �H�T$�L$ W���ĉ�T$8�H�L$<�P�H���J� �����   ;|$������L$(�T$R�T$0���ĉ�L$D�P�T$H�H�͉P�� ��u���_^][�L$(3���B	 ��,� �L$8�D$_^][3���B	 ��,� ������U��L$�����t]f�9 tWS��P  V3���~GW3��	��$    ����L  ������P�D$P�(� ����t�����   ;�|�_^[���]� ��_^[]� �U��L$�����taf�9 t[S���  V3���~KW3��	��$    �����  ���"����� P�D$P�� ����t����p;�|�_^[���]� ��_^[]� �������������Q�L$��SU�l$VWt�    �D$���  3����D$��   3�����$    �d$ �L$ �T$���  �D�;�tN��tVPVh��U�v �L$4���|$ tW��wt ���� h��U�O ����� �L$ ��t���PU���҅�t$���ø  ;t$�y���_^]3�[Y�_^]���[Y�_^]�   [Y��������������Q�L$��SU�l$VWt�    �D$��   3����D$��   3�����$    �d$ �L$ �T$���  �D�;�tN��tVPVh�U� �L$4���|$ tP��wt ���� h��U�_ ����� �L$ ��t���PU���҅�t���� ;t$|�_^]3�[Y�_^]���[Y�_^]�   [Y�����Q�L$��SU�l$VWt�    �D$��  3����D$��   3�����$    �d$ �L$ �T$��  �D �;�tN��tVPVh �U� �L$4���|$ tW��w t ���
 h��U� �����5 �L$ ��t���PU���҅�t$����  ;t$�y���_^]3�[Y�_^]���[Y�_^]�   [Y��������������Q�L$��SU�l$VWt�    �D$��   3����D$��   3�����$    �d$ �L$ �T$��  �D�;�tN��tVPVhT�U� �L$4���|$ tW��wt ��� h��U� �����E �L$ ��t���PU���҅�t$�����   ;t$�y���_^]3�[Y�_^]���[Y�_^]�   [Y��������������Q�L$��SU�l$VWt�    �D$��@  3����D$��   3�����$    �d$ �L$ �T$��<  �D�;�tN��tVPVh��U��  �L$4���|$ tP��wt ���*  h��U�  �����U  �L$ ��t���PU���҅�t����8;t$|�_^]3�[Y�_^]���[Y�_^]�   [Y�����SU�l$W�} 3�;��\$|�D$;��  |};��D$   t�L$�T$QRV�  Wh,�V�  ��8\$ t:�L$���  ��|;��  |
3�;��  }���   �E t h �V��� ����th�&V�� ���}$���|�D$;��  |]�D$��t�L$�T$QRV�� Wh��V�z� ���|$  t�����E$����t h �V�W� ����th�&V�E� ���}(���|�D$;��  |]�D$��t�L$�T$QRV�� WhؽV�	� ���|$  t�����E(����t h �V��� ����th�&V��� ����~
�D$$��t3�9D$_��][����	Ã�U3�;�VW���l$t�+�D$��0  ;ŉD$��   �l$���L$��,  |$�G;�tJ��tUPUhp�V�Y� ���|$  ��   ���ot���� h��V�2� ������� ��t��T$ �L$SRUhP����   PQ��������t�|$ u�D$	   ��BV���Ѕ�u9D$u�D$   �D$�  ��;l$�=����D$_^]���_^���]�����������Q�D$��SU�l$VWt�     �D$���  3����D$��   3ۋL$���  ���l�  ;�tV��tW���\�  PWh��U�?� ���|$ t\W���M�  ��t���� h��U�� ������� �D$ ��t� ��BU���Ѕ�t$���Ø   ;|$�r���_^]3�[Y�_^]���[Y�_^]�   [Y������Q�D$��SU�l$VWt�     �D$���  3����D$��   3ۋL$���  ����� ;�tV��tW����� PWh�U�_� ���|$ tYW���F ��t����� h��U�7� ������� �D$ ��t� ��BU���Ѕ�t!����0;|$�u���_^]3�[Y�_^]���[Y�_^]�
   [Y���������j�hHod�    P��SUW�  3�P�D$(d�    �l$@3�;�\$t�] �D$8���  ;ˉL$$u9�`  9�0  ~�D$   ;���  �\$ �	��l$@�D$8���  |$ ���� ;�t]��tS���� PSh��V�:� ���|$< t2S����D ��t���� h��V�� ������� ��t�E ��D$�������������  ���tf�}  ��   ��tSh��V��� ���|$< ��   �L$���  �L$8��@$�T$R�D$4    �ЍL$�/�  P�������t����� h��V�q� �����'� �D$@��t� ����������  �L$���D$0������  ��|$ u�D$   U�t���������   ��tSh`�V�	� ���|$< ��   �L$�"�  �L$8��R$�D$P�D$4   �ҍL$�q�  P���Y����t���>� h��V�� �����i� �D$@��t� ���W�����0�  �L$���D$0�������  ��|$ u�D$   �L$8��P U��;���   ��tPSh �V�G� ���|$< ��   �L$�`�  �L$8��@$�T$R�D$4   �ЍL$��  P�������t���|� h��V��� ������ �D$@��t� �L$�D$0������  �|$ u��BV���Ѕ�u�D$   �D$ p��;\$$�,����D$�L$(d�    Y_][��$Ã|$ ���������������̃�H�  3ĉD$D�D$XSU�l$TV�t$h3�W�|$`;��|$$�D$(�L$ �T$,�\$�\$�\$t��腣 �M;ˉL$��  3��d$ �E�\8�M�Qh`/�i���������   �D$��t�T$ SRV��� ���|$d �   �d/�`/�h/�L$4�D$0�l/�L$0Q�T$<�D$@�;������tH�T$0R�������u7�E�L$0�D$ǅ���T$4�P�L$8�H�T$<�Pt h �V�O� ����th�&V�=� ������;\$�����L$���|$$��  �U��t*�E��~#�j��t��~hjjPR诩 �L$ �����E��T$@�P�T$D�P�T$H�P�@�T$L�D$P�4  ����   �L$ �M�<Wh`/����������   �T$@RW�����������   �D$��t�G�L$P�T$,PQRV�_� ���|$d �   �d/�`/�h/�L$4�D$0�l/�L$0Q�T$<�D$@��������tH�T$0R�������u7�E�L$0�D$Å���T$4�P�L$8�H�T$<�PtDh �V��� ����t2h�&V��� ���"��O�W�D$@�G�L$D�O�T$H�D$L�L$P���l$ ������L$�|$$��tKQ���
� �|$��~;3��U�L2�2�j Q���̉�P�Q�P�@�Q�A�L$<�?� ����uǋD$(��t#�L$�T$��D$�_^][�L$D3���1	 ��HËL$�T$_^��L$L][3���1	 ��H���������������V��~ �|�t%�F��tj P����F    �F    �F    ^�����������j�hxod�    P��@�  3ĉD$<SUVW�  3�P�D$Td�    �D$d�D$(��P  3�3�;ǉL$4�T$ �|$,�D$<�=  �|$$�D$(��L  |$$����Y��������  V�i�������u�D$ ��t2VUh��P� �L$(��BV��;�t�L$ ��tPUhP�Q��� ��2ۀ|$h ��   �L$���  �t$(��R�D$P���D$`    �ҍL$�?�  P���������tP�6�L$���$�  �L$(P��Ѓ��u4�L$��  P�������D$4��t� �D$ ��th��P�G� ����L$�D$\������  ��u�|$, u�D$,   �D$$�   ��;l$<�����3�3�9|$<�l$��  �t$(�|$8��L  \$8�D$9{�\$0�|$$�  �|$�CD$��(�R���̉)�h�i�h�@�i�A���҅�}]�t$ ��t�D$$�L$PQh�V�� ���|$h ��   �S�B�KW�ЋD$4��t� ����  h��V�G� ���o  �L$(�4@���\  �N��<����t�t$ ��t��T$$�D$RPh��넃~ um�t$ ��t�L$$�T$QRh`�V��� ���|$h t4�C�P�KW�ҋD$4��t� ����   ��h��P�� ����   ���D$�D$ ��   �N��B(��=   �
  �NQ�H����������   �\$(�3�L$0�T$@R����������̉�P�Q�P�@�Q��AU���҅���   �t$ ��t�D$$�L$PQh�V�� ���|$h tk�L$0�Q�B��W�ЋD$4��t� ��t��h��Q��� ���\$0�D$$;{�t$(������l$3�9{F�D$ ;�tEUh�P�� ��3��2���D$�D$ �D$,����뭃��D$룃��D$띀|$ u9|$,u�D$,   �D$8�   ��;l$<�l$�P����D$,�L$Td�    Y_^][�L$<3��
-	 ��L������������̃�SUV���D$��`  3�3�;ÉD$��   �\$W���$    �L$��\  |$� u���   t^Sh�V�� ���M�O��Bj �Ѕ�u=���ht6Sh��V�� ������ ����� �O��BV�Ћ��,� ���%� �L$$�T$ �D$QRSh����WP���������u��t��D$�   ��;\$�E���_^��][��������������V��~ ���t%�F��tj P�ĭ�F    �F    �F    ^�����������V��F�V;�u=���Ɂ�   v��|�nff ;�}�������   ��;�}P���6����N���N��3���A�A�A�A�N�F�����N��^�������V��~ ���t%�F��tj P����F    �F    �F    �D$t	V�_�������^� ������V��~ �|�t%�F��tj P����F    �F    �F    �D$t	V��������^� ������V��~ ���t%�F��tj P�ĭ�F    �F    �F    �D$t	V��������^� ������S�\$��UVW��}P3�9nt<�~��x#��i�X  �N��P�U�҃���X  ;�}�N��PUQ���҉n_�n�n^][� �F;�}y�N��PSQ����3�;FtU�N��+�i�X  i�X  WR�Q�V.	 �F��;�}$����i�X  +�F�P���������X  ��u�_�^^][� _�V�V^][� ~X���;�|)��+�i�X  ����N�9�B�j �Ё�X  ��u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� S�\$��UVW��}P3�9nt<�~��x#��i۸  �N��P�U�҃���  ;�}�N��PUQ���҉n_�n�n^][� �F;�}y�N��PSQ����3�;FtU�N��+�iɸ  i��  WR�Q�-	 �F��;�}$����i��  +�F�P��������Ǹ  ��u�_�^^][� _�V�V^][� ~X���;�|)��+�i��  ����N�9�B�j �Ё�  ��u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� S�\$��UVW��}K3�9nt7�~��x����N��P�U�҃���0;�}�N��PUQ���҉n_�n�n^][� �F;�}{�N��PSQ����3�;ǉFtW�V��+ʍI�R��Q���WR��+	 �F��;�}&�<@����+荤$    �F�P��������0��u�_�^^][� �~�~_^][� ~S���;�|$�<@+�������N�9�B�j �Ѓ�0��u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� ��������S�\$��UVW��}J3�9nt6�~��x�����N��P�U�҃��� ;�}�N��PUQ���҉n_�n�n^][� �F;�}m�N��PSQ����3�;FtI�N��+���W��R�Q�*	 �F��;�}������+�F�P�������� ��u�_�^^][� _�V�V^][� ~R���;�|#��+�������N�9�B�j �Ѓ� ��u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� ��������S�\$��UVW��}P3�9nt<�~��x#��i�  �N��P�U�҃���  ;�}�N��PUQ���҉n_�n�n^][� �F;�}y�N��PSQ����3�;FtU�N��+�i�  i�  WR�Q�f)	 �F��;�}$����i�  +�F�P���c�����  ��u�_�^^][� _�V�V^][� ~X���;�|)��+�i�  ����N�9�B�j �Ё�  ��u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� S�\$��UVW��}P3�9nt<�~��x#��i��   �N��P�U�҃����   ;�}�N��PUQ���҉n_�n�n^][� �F;�}y�N��PSQ����3�;FtU�N��+�i��   i��   WR�Q�&(	 �F��;�}$����i��   +�F�P����������   ��u�_�^^][� _�V�V^][� ~X���;�|)��+�i��   ����N�9�B�j �Ё��   ��u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� S�\$��UVW��}W3�9ntC�~��x*��    +���ۍI �N��P�U�҃���8;�}�N��PUQ���҉n_�n�n^][� �F;���   �N��PSQ����3�;ǉFtg�V��+ʍ,�    +����    �U+ʍ�WR��&	 �F��;�})�<�    +������+萋F�P���c�����8��u�_�^^][� �~�~_^][� ~a���;�|2�<�    +���+��������I �N�9�B�j �Ѓ�8��u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� ����������S�\$��UVW��}P3�9nt<�~��x#��i��   �N��P�U�҃����   ;�}�N��PUQ���҉n_�n�n^][� �F;�}y�N��PSQ����3�;FtU�N��+�i��   i��   WR�Q�v%	 �F��;�}$����i��   +�F�P���c������   ��u�_�^^][� _�V�V^][� ~X���;�|)��+�i��   ����N�9�B�j �Ё��   ��u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� V��~ ��t%�F��tj P���F    �F    �F    ^�����������V��~ �4�t%�F��tj P�@��F    �F    �F    ^�����������V��~ ��t%�F��tj P���F    �F    �F    �D$t	V���������^� ������V��~ �4�t%�F��tj P�@��F    �F    �F    �D$t	V��������^� ������SW�|$����~mU�l$��|cV�t$��|Y;�tU�C�/;�K;�G�K�>;�~�;�}��P���f���C����+��ҋ���+�R������R+΍�R�#	 ��^]_[� ��U�l$V��;�t[�ES3�;��^[��^]� 9F}P����9^t�E;ÉF~�W3����E�N�P����������X  ;^|�_[��^]� ��^]� ��j�h�od�    PQSVW�  3�P�D$d�    ���|$���   3�9^�D$   ��t�F;�tSP�����^�^�^9��   ���   �D$��t�F;�tSP�����^�^�^9��   ���   �D$��t�F;�tSP�����^�^�^9��   �wt�D$��t�F;�tSP�����^�^�^9_p�wd�D$��t�F;�tSP�����^�^�^9_`�wT�\$��t�F;�tSP�����^�^�^9_P�wD�D$������t�F;�tSP�����^�^�^�L$d�    Y_^[������������������j�hpd�    P��@  �x)	 �  3ĉ�$�@  SUVW�  3�P��$�@  d�    ��$�@  ��$�@  3�;Ë���   hD�P�l� ����;�tpVj�L$�'� j�L$��$�@  襡 j�L$�ʡ j�L$�� ��$�@  ��$�@  UPQ�T$ R������V���� ���L$Ǆ$�@  ������ �Ë�$�@  d�    Y_^][��$�@  3��z	 �ļ@  � �������j�hXpd�    P��SUV�  3�P�D$$d�    ��`  ���  3�3�襉 ;��  S�L$�D$���l$�l$ �l$$�϶��;݉l$,~>�\$�I ��\  �L$��/����N��V�P�N�H�V���   �l$�Pu�3�D$<�L$8�T$4PQR���  P�D$$P�x��H��?�������;�tP�|$4 tI;�~E3����$    �L$��\  �
�H�I���L)�(�)�h�i�h�i�@�����Au�3�9l$ �D$,�����D$��t�D$;�tUP�L$����ƋL$$d�    Y^][�� ��������j�h�pd�    P��D�  3ĉD$@UVW�  3�P�D$Td�    �D$h����0  3�D$ 3�;��|$�l$�t$�#  V�L$(�D$(���l$,�l$0�l$4�I������l$\�(  �l$���$    ��,  D$���   �pWV�V���������   �D$��tUh0�S�F� ���|$d t]�D$ ��t� Vh`/薫������t��W�G��O�V�F�N���F�N��V�G�O�W��t h �S��� ����th�&S��� ��Vh`/�2��������L$$t��������W�P�O�H�W���������V�P�N�H�V�D$�  �|$��;l$�P������t$�D$ �L$dSPQ�T$0j R������������D$�D$to�|$d th��~d3ҋD$(�,��Ai��  �,  �����h�i�h�i�h�I�H�H���   �H���   �H���   �H���   u��t$�D$3�;��l$��  ���  �T$4��,  �D$8P��D$<�����N�V���ĉ�N�P�V�H�L$H�P�v� ����  �D$��t�D$8�L$PQh��S�P� ���|$d �G  �L$<�٪ �`/�h/3��D$<�D$@�D$D�D$H�D$L�d/�D$@�T$<�l/�D$<P�L$H�T$L�D$P��������������   �L$<Qh`/�@���������   �T$<�L$@P���ĉ�T$X�H�L$\�P�H�L$H蛑 ����   �L$(��t;�D$,��~3hPjjPQ�T$LR�b5	 ����t+D$(�ȸgfff���������yU�D$ ��t� �ۋD$<�L$@�T$D�|$H�F���   �N���   �V���   �~���   t&h �S�� �|$ ����th�&S��� ����|$�D$���Ő  ;D$�D$�����D$�|$0 �D$\�����D$$��t�L$(��tj Q�L$,����D$�L$Td�    Y_^]�L$@3��d	 ��P�������j�h�pd�    P��SUV�  3�P�D$$d�    ��P  ���  3�3�蕃 ;��  S�L$�D$���l$�l$ �l$$述��;݉l$,~>�\$�I ��L  �L$������N��V�P�N �H�V$���   �l$�Pu�3�D$<�L$8�T$4PQR���  P�D$$P����h��/�������;�tP�|$4 tI;�~E3����$    �L$��L  �
�Hi��   �L)�(�)�h�i�h�i�@�����Au�3�9l$ �D$,�����D$��t�D$;�tUP�L$����ƋL$$d�    Y^][�� ��������j�h�pd�    P��SUV�  3�P�D$$d�    ���  ���  3�3��%� ;��  S�L$�D$���l$�l$ �l$$�O���;݉l$,~>�\$�I ���  �L$������N��V�P�N�H�V�Ÿ  �l$�Pu�3�D$<�L$8�T$4PQR���  P�D$$P��������������;�tP�|$4 tI;�~E3����$    �L$���  �
�Hiɸ  �L)�(�)�h�i�h�i�@�����Au�3�9l$ �D$,�����D$��t�D$;�tUP�L$����ƋL$$d�    Y^][�� ��������j�hqd�    P��SUV�  3�P�D$$d�    ���  ���  3�3�赀 ;��  S�L$�D$���l$�l$ �l$$�߭��;݉l$,~>�\$�I ���  �L$��?����N��V�P�N�H�V�Ř   �l$�Pu�3�D$<�L$8�T$4PQR���  P�D$$P�D����O�������;�tP�|$4 tI;�~E3����$    �L$���  �
�Hiɘ   �L)�(�)�h�i�h�i�@�����Au�3�9l$ �D$,�����D$��t�D$;�tUP�L$����ƋL$$d�    Y^][�� ��������j ����������̃�SU�l$W��SV��U�D$    �r���������   ~�L$�ɉD$t�D$P�D$   臶��VU������������   ~�L$D$��t�T$R�D$   �S���SVU����������   ~�L$D$��t�D$P�D$   � ���SVU�X�������|S~�L$D$��t�T$R�D$   ����SVU��������|$~�L$D$��t�D$P�D$   �µ���D$_][����������j ���������UW��3�9o��t;V�w��x S�v���O��P�U�҃���0;�}�[�O��PUQ���҉o^�o�o_]�������������t���������̋D$SU�@V�t$��PV���&���������t)��t%;�t!W3�9{~����B���Ѓ���0;{|��_^][� ��������������V��V2���tQ�N��~JW�|$��t@��~9Wj0QR资 3���9~~%S3����    �F���B�Ѓ���0;~|�[�_^� ���������������V��V2���tQ�N��~JW�|$��t@��~9Wj0QR�5� 3���9~~%S3����    �F���B�Ѓ���0;~|�[�_^� ���������������SUVW�|$����t�    �D$ �\$P�D$ S�t$ �D$     ���������t�L$����  �t$V�T$RSU�D$0�D$(    ���������t�L$����  V�T$RSU�D$(    ��������t�L$���t  V�T$RSU�D$(    ��������t�L$���J  �T$RSU�D$$    �n�������t�L$���!  V�T$RSU�D$(    �4�������t�L$����   V�T$RSU�D$(    ���������t�L$����   V�T$RSU�D$(    ��������t�L$����   SU�ƍ\$ �D$     ���������t�T$��|}�ދt$S�D$PVU�D$(    �J�������t�L$��|QVU�ӍL$ �D$     ��������t�T$��|+�D$PVU���D$$    ��������t�L$��|�D$ _^][� �UW��3�9o�0�t:V�w��xS��k�p�O��P�U�҃���p;�}�[�O��PUQ���҉o^�o�o_]������������������������̋D$k�pSUV�t$PV���Y���������t)��t%;�t!W3�9{~����B���Ѓ���p;{|��_^][� �V��V2���tQ�N��~JW�|$��t@��~9WjpQR��� 3���9~~%S3����    �F���B�Ѓ���p;~|�[�_^� ���������������V��V2���tQ�N��~JW�|$��t@��~9WjpQR�u� 3���9~~%S3����    �F���B�Ѓ���p;~|�[�_^� ���������������UW��3�9o�D�t:V�w��xS�����O��P�U�҃��� ;�}�[�O��PUQ���҉o^�o�o_]������������������������̋D$SUV�t$��PV������������t)��t%;�t!W3�9{~����B���Ѓ��� ;{|��_^][� �V��V2���tQ�N��~JW�|$��t@��~9Wj QR�U 3���9~~%S3����    �F���B�Ѓ��� ;~|�[�_^� ���������������V��V2���tQ�N��~JW�|$��t@��~9Wj QR��~ 3���9~~%S3����    �F���B�Ѓ��� ;~|�[�_^� ���������������j �X��S������j �l��������j ����������j ����������VW�|$����|o;~}j�N����j<+Ǎ�j R��	 �F��+ǃ�P�OQW���0����F����+ЋFj<�L��j Q��	 �F����+ЋF�L�ă�Q�������F�_^� V��j ���������D$t	V�C�������^� ����������V��������D$t	V��������^� ��V���t�������D$t	V���������^� ������������V���x����D$t	V���������^� ��V������R����D$t	V��������^� ������������V��������D$t	V�{�������^� ��V����������D$t	V�U�������^� ������������V��j �l������D$t	V�#�������^� ����������V��j ����0����D$t	V���������^� ����������SVW�|$����}@3�9^��   �~��x�F����l ��y���F�RSP����_�^�^�^^[� �F;�}[�N��PWQ����3�;ÉF��   �N��+����R��SP�
	 �^��;�}�N��R���������;�|�~_^[� ~H�X�;�|��$    �F���El ��;�}�9~~�~��F�RWP�Ή~��3�;ÉFu�^�^_^[� j�hKqd�    P��  �  3ĉ�$�  SUVW�  3�P��$�  d�    ��$�  ��F�n;���   ��iɸ  ��   v��|��� ;�}�ȍ<����   ~�< �F��tz��+ȸ� O	���������xc;�}_�L$�A�  S�L$Ǆ$�      ��}  9~}W�������F��iɸ  N�T$��R�F�}  �L$Ǆ$�  �����}  �&;�}W���_����F��iɸ  N��S�F�e}  ��$�  d�    Y_^][��$�  3��.	 ���  � ����������̋D$i��  SUV�t$PV�������������t,��t(;�t$W3�9{~����B���Ѓ��Ƹ  ;{|��_^][� �����������V��V2���tT�N��~MW�|$��tC��~<Wh�  QR�ry 3���9~~%S3���I �F���B�Ѓ��ø  ;~|�[�_^� ������������V��V2���tT�N��~MW�|$��tC��~<Wh�  QR��x 3���9~~%S3���I �F���B�Ѓ��ø  ;~|�[�_^� �����������̋D$i��   SUV�t$PV������������t,��t(;�t$W3�9{~����B���Ѓ��Ƙ   ;{|��_^][� �����������V��V2���tT�N��~MW�|$��tC��~<Wh�   QR�2x 3���9~~%S3���I �F���B�Ѓ��Ø   ;~|�[�_^� ������������V��V2���tT�N��~MW�|$��tC��~<Wh�   QR�w 3���9~~%S3���I �F���B�Ѓ��Ø   ;~|�[�_^� ������������V��j ���s���D$t	V���������^� ����������j�h�qd�    P��4�  3ĉD$0SUVW�  3�P�D$Hd�    �\$X���G�o;���   �@����   v��|���* ;�}�ȍ4����   ~�4 �G��tr��+ȸ���*���������x[;�}W�L$� S�L$�D$T    �=���9w}V��������G�@��O�T$��R�G�����L$�D$P������ �_;�}V�������G�4@��w��S�ΉG�{����C�F�K�N�S�V�C�F�K�S�NR�N�1�  �F �P�N �� S�ҋL$Hd�    Y_^][�L$03�� 	 ��@� �j�h�qd�    P��$�  3ĉD$ SVW�  3�P�D$4d�    �\$D���G�W;���   ������   v��|� @ ;�}�ȍ4����   ~�4 �O��tc��+���xZ;�}V�L$��s S�L$�D$@    �ݝ��9w}V��������G����O�T$��R�G赝���L$�D$<�����$t �S;�}V�������G����w��S�ΉG�����CP�N���  �K�C�N��N��P�Q�P�Q�@�A�L$4d�    Y_^[�L$ 3��� ��0� ���������������j�h�qd�    P��  �  3ĉ�$  SUVW�  3�P��$0  d�    ��$@  ��F�n;���   ��i�  ��   v��|�}P ;�}�ȍ<����   ~�< �F��t|��+ȸ������������xc;�}_�L$�_� S�L$Ǆ$<      誜��9~}W���m����F��i�  N�T$��R�F�����L$Ǆ$8  �����;� �&;�}W���-����F��i�  N��S�F�C�����$0  d�    Y_^][��$  3��L� ��(  � ��������̋D$i�  SUV�t$PV������������t,��t(;�t$W3�9{~����B���Ѓ���  ;{|��_^][� �����������V��V2���tT�N��~MW�|$��tC��~<Wh  QR�r 3���9~~%S3���I �F���B�Ѓ���  ;~|�[�_^� ������������V��V2���tT�N��~MW�|$��tC��~<Wh  QR�r 3���9~~%S3���I �F���B�Ѓ���  ;~|�[�_^� ������������V��j �X������D$t	V�C�������^� ����������j�h+rd�    P���   �  3ĉ�$�   SUVW�  3�P��$�   d�    ��$�   ��F�n;���   ��i��   ��   v��|�x=
 ;�}�ȍ<����   ~�< �F��tz��+ȸ��Q���������xc;�}_�L$�� S�L$Ǆ$�       �|���9~}W��������F��i��   N�T$��R�F�Q����L$Ǆ$�   ������ �&;�}W�������F��i��   N��S�F������$�   d�    Y_^][��$�   3��~� ���   � ����������̋D$i��   SUV�t$PV���6���������t,��t(;�t$W3�9{~����B���Ѓ����   ;{|��_^][� ����������̋D$S�ٍ�    +��U�V�t$�QV�����������t+��t';�t#W3�9{~������B���Ѓ���8;{|��_^][� ���V��V2���tQ�N��~JW�|$��t@��~9Wj8QR�eo 3���9~~%S3����    �F���B�Ѓ���8;~|�[�_^� ���������������V��V2���tQ�N��~JW�|$��t@��~9Wj8QR��n 3���9~~%S3����    �F���B�Ѓ���8;~|�[�_^� ���������������V��j ���������D$t	V��������^� ����������j�hkrd�    P���   �  3ĉ�$�   SUVW�  3�P��$�   d�    ��$�   ��F�n;���   ��i��   ��   v��|�x=
 ;�}�ȍ<����   ~�< �F��tz��+ȸ��Q���������xc;�}_�L$�Q���S�L$Ǆ$�       ����9~}W���_����F��i��   N�T$��R�F�����L$Ǆ$�   �����-����&;�}W�������F��i��   N��S�F赟����$�   d�    Y_^][��$�   3��N� ���   � �����������V��V2���tT�N��~MW�|$��tC��~<Wh�   QR��l 3���9~~%S3���I �F���B�Ѓ����   ;~|�[�_^� ������������SUVW�|$����}U3�9n�  �~��x$������    �F�L�d� ����0;�}��F�RUP����_�n�n�n^][� �F;�}k�N��PWQ����3�;ŉF��   �V��+ʍI�R��Q���UR��� �F��;�}�@����+�F�P��������0��u�~_^][� ~T���;�|%�@+�������d$ �N�L褉 ��0��u�9~~�~��F�RWP�Ή~��3�;ŉFu�n�n_^][� �������������j�h�rd�    P��SUVW�  3�P�D$d�    �ى\$3��K�{�{�s����K�[ ���   �Q ��p  3�;�~%�d$ ��l  ��;�t	��Bj�Ѓ�;�p  |ߋ�l  ;�t��t  ;�~��QWP�� ��3�9��  ~#�����  ��;�t	��Pj�҃�;��  |ߋ��  ;Ǎ��  t�N;�~��QWP�<� ��9~t�F;�t�WP�B���Љ~�~�~9��  ���  tK�u��x1��i��  �D$��$    �ML$W��B�Ёl$�  ��;�}�U �E�RWP���҉}���  �}�}9~tC�n��x*��i��   �D$�NL$W��P�ҁl$�   ��;�}�N��PWQ���҉~�~�~9��  ���  t<�n��x�\m ���N��P�W�҃���0;�}�N��PWQ���ҋ\$�~�~�~9��  ���  tD�n��x+��k�p�D$��$    �NL$W��P�҃l$p��;�}�N��PWQ���҉~�~�~9��  ���  t=�n��x$�����D$�NL$W��P�҃l$ ��;�}�N��PWQ���҉~�~�~9�  ��  tC�n��x*��i�  �D$�NL$W��P�ҁl$  ��;�}�N��PWQ���҉~�~�~9�  ��  tH�n��x+��i��   ���    �N��P�W�҃����   ;�}�N��PWQ���ҋ\$�~��(  �~�~9}te�}��x@��iې  �u�t$���   �D$$   ������D$$�����M  ����  ��}ȋM�E �Pj Q���ҋ\$�E    3��}�}9�<  ��8  tE�u��x'��    +���ۋM��P�W�҃���8;�}�M�E �PWQ���ҋ\$�}��H  �}�}9~t@�n��x#��i��   �N��P�W�҃����   ;�}�N��PWQ���ҋ\$�~�~�~9�\  ��   ��d  ����   �Dm ���D$����D$��\  ��t$���   ;��D$$   t 98v� ����   98wP����������   9��   u�N;�t�> t	��Pj�ҍN�~� �D$$���������l$�   ��;��x�����\  ��X  �P��X  WQ���҉~��h  ��`  ��d  9~t�F;�t�WP�B���Љ~�~�~9�|  ��x  tH�u��x.�v���D$���    �M�T$�L
萃 �l$0��;�}�M�E �PWQ���҉}�}�}���  ���  ���  ��] ���  ��] ���  ��] ���  ��] ���  �j �L$d�    Y_^][��������VW�|$W���R����G�F�O�N�W�V�G�F�O�W�NR�N��  �G P�N ���  �O$�N$�W(�V(�G,�F,�O0�N0�W4�V4�G8�F8�G@�^@�GH�^H�GP�^P�GX�^X�O`�N`�Wa�Va�Gb�Fb�Oc�Nc�Gd�Nd;�tP�����Vt�R�Nt�GtP�ҋ��   ���   ���   �P���   �H���   �P_���   ��^� ��̃�SUVW���L$(�I3����D$�L$�  ����+����D$ ��D$ �T$(�j�]4�ۍE4�D$|/�G0�O�WPQ�wdR��芘����;؉D$t�L$�D$��� �����]8��|,�W0�O�GRPQ�wd���N�����;؉D$t�D$�E8��E8�����T$������   ;G��   �i��   ���  �u�DVP����������   V�D$�����U�������uI��L$Q�N���ĉ�V�H�N�P�H����  �!h ��t�D$��|;G}�T$��   �D$��iɘ   ���  �D���P�V�H�N�P�V�\�uVh`/�7������t�D$� �����;�L$�Q�N���ĉ�V�H�N�P�H����  �g ��u
�T$������E8����]8��   ;G��   �i��   ���  �u �DVP�~��������   V�D$�����,�������uB��L$Q�N���ĉ�V�H�N�P�H����  ��f ��t�D$��|	;G}��t��iҘ   ���  �D
���H�N�P�V�@�F�H�u Vh`/�~������u-��VS���ĉ�N�P�V�H����  �P�yf ��u������D$�8 }�; }�L$Q�L$,������D$�l$ <�����D$�����D$_^][��� �������������S�\$UVW�sV��3���������tV�������   �G4�W�KDP�GR�wtP�L$ �j�����9D$t�CD���W0�G�K0R�WP�wdR�L$ �?�����9D$t�C0����4S���5���_^�][� ������������j�h�rd�    P��SUVW�  3�P�D$(d�    �ًl$8�uV�D$    �B�������tV��������D$   �C(�K�S�} PQ�sDR��蠔����;�t�D$�E �C4�K�S�}$PQ�stR���w�����;�t�D$�E$�C0�K�S�}(PQ�sdR���N�����;�t�D$�E(���������  3��D$�$�D$�D$ �D$$�D$0�D$P���y���|$ ���3�;��}   �sT��I �L$�,��S,�K�CRPQ���Փ������}8��|?�D$ ;�}7+ǃ�P�WRW�L$$������D$ �L$���D$ ��    �;�t�T$���D$��y��l$83����$��3�9t$ ~�D$��Q��������;|$ |�9t$$�D$0�����D$�$t �D$;�tVP�L$ ��$�t$�t$$�t$ ��,U���#���D$�L$(d�    Y_^][�� � ���������SV��3�9^�h�t1W�~��x��    �F���N ��y���F�RSP���҉^_�^�^^[������j�hsd�    P��H�  3ĉD$DSUVW�  3�P�D$\d�    �D$p�T$x�t$l���L$t�L$L�D$H�D$|�L$HQ�T$T�D$X��������t3��l  �F�N�V�D$<�D$8�L$@�T$8�VP�L$LQ�T$L�e�������u
�   �0  �L$8��R���ĉ�L$L�H�L$P�H�L$T�H���҃��u���  i��   �L  3�h   3�U�L$�؉t$0�D$4��l$ �l$$�l$(�@�;ŉD$t7�L$ ��   }�   +���R��UP�[� �D$$���T$�D$    �
3҉l$ �T$�K;͉l$d�l$$��   �C�4(��RŃ��̉1�p�q�p�@�q�A���҅�|Z�4@���\  �~ tH�N��P(��=   u7�FP���������D$0t#��P�L$LQ���������L$t:�T$0R聯���D$$����;C�D$$�a����T$�D$�t$(3�   �\$,�%�D$d����������   �  ���$    ��t$(;��E  ��;ʉT$(�L$4�  ����3�;���   �Y��R�A���̉�X�Y�X�@�Y�A����;���   i��   �L  �l$$��9k��   �C�4(��RŃ��̉1�p�q�p�@�q�A���҅�|^�4@���\  �~ tL�N��P(��=   u;�FP辂�������D$0t'��P�L$LQ�����������   �T$0R�L$�,����D$$����;C�D$$�]����t$4�D$��;t$(�t$4������T$�\$,��3���  �\$,�����3Ɂ��  ���D$d�����D$4������9l$ ��t;�tUP�L$�@��ƋL$\d�    Y_^][�L$D3��� ��T� �|$  �D$d�����D$4�t�D$��tj P�L$�@��D$,��UV��3�9n���t<W�~��x!S��iې  �N��z������  ;�}�[�N��PUQ���҉n_�n�n^]�����������UW��3�9o���t:V�w��xS�v���O��e|�������   ;�}�[�O��PUQ���҉o^�o�o_]�������������UW��3�9o�̭t9V�w��xS�v���G�L�v ����0;�}�[��G�RUP���҉o^�o�o_]��������������V���X����D$t	V���������^� ��V�������D$t	V�ۨ������^� ��V��������D$t	V軨������^� ��V���8����D$t	V蛨������^� ��j�h;sd�    P��   �  3ĉ�$�   SUVW�  3�P��$�   d�    ��$�   ��F�n;���   ��iɘ   ��   v��|�Ky ;�}�ȍ<����   ~�< �F��tz��+ȸ��k���������xc;�}_�L$�1�  S�L$Ǆ$�       �,���9~}W���S���F��iɘ   N�T$��R�F�����L$Ǆ$�   ����譐  �&;�}W���?S���F��iɘ   N��S�F�������$�   d�    Y_^][��$�   3���� �Ĩ   � �����������V��F�V;�uP�@����   v��|���* ;�}�������   ��;�}BP�������N�I��F���N^Í@�F���L�1t �F�@��NQ���M����N�I��F���N^����������j�h�td�    PQSUVW�  3�P�D$d�    ��t$3��^���(��~�~�-|���n�͉|$ �_� ���   �D$ ��> ǆ�  |����  ���  ���  ���  ���  ���  ǆ�  �����  ���  ���  ǆ�  �����  ���  ���  ǆ�  t����  ���  ���  ǆ�  �����  ��   ��  ǆ�  ����  ��  ��  ǆ  ����  ��   ��$  ǆ  ��ǆ(  ����,  ��0  ��4  ��<  ��@  ��D  ǆ8   ���L  ��P  ��T  ǆH  �ǆX  ����\  ��`  ��d  ǆh  ����l  ��p  ��t  ǆx  ̭��|  ���  ���  ���  �D$ �X ���  �D$ �wX ���  �D$ �gX ���  �D$ �WX ���  �D$ ���  ���  �X ���D$ ��}������� ���   �-: �ƋL$d�    Y_^][����������j�h�ud�    PQSVW�  3�P�D$d�    ��t$�(��D$   ��������  �D$�X ���  �D$�#X ���  �D$�X ���  �D$�X ���  �D$��W ��x  �D$������h  3�9_�D$���t�G;�tSP���ĭ�_�_�_��X  �D$�a�����H  S�D$ ����J�����8  S�D$ ����ù����(  �D$
�������  S�D$ 	�l��\�����  S�D$ �X��������  �D$�����������  �D$����9������  �D$�t��S������  S�D$ ���,N�����  S�D$ �������9��  ���  �D$�|�t�G;�tSP������_�_�_���   �D$�b< �N�\$�� �N�D$�����f{���L$d�    Y_^[������SUV�t$3��W����   ��P(���҃�@��   =   tD=   ��   V�5 ��������   ����. ��V���t���;�tqP����. _^��][� V�ً ������tQ���I� �����   ��Wt	�����;������;�t+_���   �   ^��][� V��������t
P��������_^��][� �����̃�SUVW����W(���  �GR�WP3�wDR�l$��������|;G|3����k�p���  ����  ��j�����u"����  j��%�������  j ��d�������  �W(3�9��  ~*3ۋ���  �P������������p;��  |܉l$���    �D$    ��   3� ���  �\)l�W8�G�T$�D$��tO3��D$ �D$$���   ���\$ t7���   ��~-h &jQP�L$0Q�w� ����t���   +�����|�t���|;t$|�t$;�t���  �D$�t(l�D$������   ;�   �D$�M����l$�3�9�0  ~93ۍ�$    ���,  ��   P���y�������Ð  ;�0  |ԉl$�3�9�`  ~P3�����\  �L.�Q���*�����V�ωD$ �+���D$�D$�����   ;�`  |��D$_^][���_^��][�������������S�\$��UVW��}|3�9~th�^��xO�,�    +����I �F�|(4 �|((�%t�G��tj P���%3��G�G�G����8��}�3���F�RWP���҉~�~�~_^][� �F;���   �N��PSQ����3�;ǉFtf�V��+ʍ,�    +����    �U+ʍ�WR�)� �F��;�}(�<�    +������+�F�P����x����8��u�_�^^][� �~�~_^][� ��   ���;�|^�,�    +���+����D$�	��$    ���N�|)4 �|)(�%t�G��tj P���%3��G�G�G��8�l$u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� ������j�hvd�    P��t�  3ĉD$pSUVW�  3�P��$�   d�    ��$�   ��F�n;���   ��k�p��   v��|�,I ;�}�ȍ<����   ~�< �F��ty��+ȸ�$I�����������x`;�}\�L$�x���S�L$Ǆ$�       �S���9~}W���VI���F��k�pN�T$��R�F�+����L$Ǆ$�   ���������#;�}W���I���F��k�pN��S�F�������$�   d�    Y_^][�L$p3��^� �Ā   � �����������U�l$V��;�tX�ES3�;��^[��^]� 9F}P�����9^t�E;ÉF~�W3����E�N�P��P������8;^|�_[��^]� ��^]� �����V���(����D$t	V�+�������^� ��j�hqvd�    P��`  �  3ĉ�$\  SUVW�  3�P��$t  d�    �����  3�3����\$~f����  ����u���  �P���  W���҃��,9xt�x���hUh`/�f������tU�Э���������;��  |��\$����  �lB ����  Q���  �E �3�9��  ~z3ۋ���  �9ht�D$�h�xWh`/�5f������tW�X������D$��Wj U���ĉ�O�P�W�H����  �P�R ����ø  ;��  |�����  ��A ����  Q���  ��D ��F ���  �^d3�F9k|�k�F9C}P���u���9n��   �l$���    ����  �C�S|$;�u=��    ��   v��|�  ;�}�������   ��;�}P�������S�K3��щD��C�ыS���C�i�G�9ot�D$�o�F��Wh`/��d������tW�������D$��Wj U���ĉ�O�P�W�H����  �P�5Q �D$�   ��;n������F ���  �^t3�F9k|�k�F9C}P���E���9n��   �D$    �d$ ����  �C�S|$;�u=��    ��   v��|�  ;�}�������   ��;�}P��������S�K3��щD��C�ыS���C�i�G�9ot�D$�o�F��Wh`/�c������tW�ت�����D$�D$0��;n�?�������  ����   �L$ �u���3��L$ ��$|  �C������R$��$�   P�ҍ�$�   �v�  P� f������uhP���$�   ��  �D$,P�|$,�J������L$ Q����  ������D$�L$ Ǆ$|  �����L�����F ���  �^D3�F9k|�k�F9C}P������9n��   �l$�I ����  �C�S|$;�u=��    ��   v��|�  ;�}�������   ��;�}P���=����S�K3��щD��C�ыS���C�i�G�9ot�D$�o�F��Wh`/�b������tW�8������D$�D$p��;n�?�����F ��   �^T3�F9k|�k�F9C}P������9n��   �D$    ������  �C�S|$;�u=��    ��   v��|�  ;�}�������   ��;�}P���=����S�K3��щD��C�ыS���C�i�G�9ot�D$�o�F��Wh`/�a������tW�8������D$�D$ ��;n�?�����   9�  ��   ��$X  ��� ��$X  ��$|  �� ��$`  ��  P�c������uhP���$d  胖  ��$|  RǄ$|      諧�������$X  P��  �C���|$��$X  Ǆ$|  �����h� ��F ��  ���   3�F9k|�k�F9C}P�������9n��   �D$    ���    ���  �C�S|$;�u=��    ��   v��|�  ;�}�������   ��;�}P�������S�K3��щD��C�ыS���C�i�G �9o t�D$�o �F��$Wh`/�e_������tW舦�����D$�D$  ��;n�<�����   9�   ��   ��$�   �� ��$�   Ǆ$|     �� ��$�   �*�  P��a������uhP���$�   �̔  ��$�   3�R��$�   ����������$�   P��  ��$   �W���|$��$�   Ǆ$|  �����L� �3��F	 ��   ���   �V 9k|�k�F 9C}P���;���9n ��   �D$    ���  �C�S|$;�u=��    ��   v��|�  ;�}�������   ��;�}P��������S�K3��щD��C�ыS���C�i�G�9ot�D$�o�F	��Wh`/�]������tW�Ҥ�����D$�D$�   ��;n �<����3�9�0  �L$��   �\$�L$����    �L$���,  D$9Ht�H�����   �xUW�5]������Wh`/��   �]������t#W�B�������W�G�M �O�U�E�M���D$��D$�  ��;�0  �D$�t����\$��F
 ��@  ���   3�N$9k�\$|�k�F$9C}P���}���9n$�&  �D$    ���<  �C�S|$;���   ��    ��   vn��|i�  ;�}����h�J\������t�U �E�M��U�G�O�W�/���Uh`/�\������������O�W�E �G�M�U�E��������   ��;�}P�������S�K3��щD��C�ыS���C�i�G;�t�D$�o�F
��Wh`/�[������tW跢�����D$�D$8��;n$���������  �Q7 ���P  Q���  �m: �3�9�P  ~m3ۋ��L  ÍxWh`/�'[������tW�J������D$��Wj U���ĉ�O�P�W�H����  �P�wG ������   ;�P  |�����  �6 ���`  Q���  ��9 �3�9�`  ~r3���I ���\  ÍxWh`/�Z������tW諡�����D$��Wj U���ĉ�O�P�W�H����  �P��F ������   ;�`  |���l$3�9�p  ~S���l  ����u��h  ��PW���҃��!�Y Sh`/��Y������tS�����������;�p  |��~ t-�NH��t&�FL��~�0&��t��~h0&jPQ��< ���~ t-�NX��t&�F\��~�0&��t��~h0&jPQ�< ���~ t-�Nh��t&�Fl��~�0&��t��~h0&jPQ�< ���~ t-�Nx��t&�F|��~�0&��t��~h0&jPQ�Y< ���~ t3���   ��t)���   ��~�0&��t��~h0&jPQ� < ���~	 t3���   ��t)���   ��~�0&��t��~h0&jPQ��; ���~
 t1�D$�H��t&�@��~�0&��t��~h0&jPQ�; ���ŋ�$t  d�    Y_^][��$\  3��� ��l  ����VW�|$W����a���G�OQ�N�F萌  �W�V�G�F�O�N�W�O$�V�G Q�N$�F �f�  ��(W�N(�
���_��^� ���j�h�vd�    PQV�  3�P�D$d�    ��t$�D$����3��N,�N0�N4�N@�F�F�F�F�F�F	�F
�F�F�F�F�F�F �F$�F(�F8�F<���ND�FH�FL�FP�D$�NT�FX�F\�F`�Nd�Fh�Fl�Fp�Nt�Fx�F|���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���D$�����ƋL$d�    Y^��� ���������j�h+wd�    P��   V�  3�P��$�   d�    �񍎈  �i2 ���  �^2 ���  �S2 ���  �H2 ���  �? �~d u�N�?� V�L$�e����L$Ǆ$�       �����L$Ǆ$�   �����m�����$�   d�    Y^���   �������j�hXwd�    P��<�  3ĉD$8SUVW�  3�P�D$Pd�    �\$`��F�n;���   ��    +���Ɂ�   v��|�Q�$ ;�}�ȍ<����   ~�< �F��tz��+ȸ�$I�����������xa;�}]�L$�3 S�L$�D$\    ����9~}W���ş���F�N��    +ЍэT$��R�F������L$�D$X������3 �*;�}W��脟���F�V��    +ȃ���S�F�����L$Pd�    Y_^][�L$83��%� ��H� �����U����j�hqxd�    P��`  �  3ĉ�$X  SVW�  3�P��$p  d�    �}�u�ى\$�|$$�D$     �D$�.����CP�KQ����� ��u��th(�V謄 ��2��\  ���+Q ��9��  t-��th�h��V�}� h�V�r� �����  �D$ �L$$�CP�� ��u��t�h��V�D� ��2���  �L$$h��V����Z������t�D$ �|$$���� ���   R�ωC�� ��u���L���h8�V�� ��2��  �L$$h �V���Z������t�D$ �|$$���B ����   �D$P���D$    ��S ��te};��t2h��V臃 �D$(����=�  �D$ �����h�V�c� ���D$ �L$Q���  軉���T$R���D$    �S ��u������ ��u���w���hx�V�� ��2���  �L$$hd�V���Y������t$���th��V�� h�V�ׂ ���D$ �L$$�6E ���~  �|$$�D$3�P�ω\$��b ����   }?����   h��V苂 �D$(����=�  �D$ �����h�V�g� ���   �L$,�6N���D$,(6�L$Q�L$0Ǆ$|      ��$ �|$�T$�Ǹ  R��菹���D$�X�G��~�Oi��  ��H����3�j P�L$4��$ �L$��t	��Bj�ЍL$,�D$    Ǆ$x  �����tU���|$$�L$Q�σ���a ���	������ұ ��u�������h �V苁 ��2��;  �L$$�N �\$��9��  tL��th��h��V�V� h�V�K� �����  ���thx�V�1� h�V�&� ���D$ �L$$�D ����  �L$$�T$3�R�\$�id ;��$  ��}s��t2h �V�ހ �D$(����=�  �D$ ����h�V躀 ��h�   ��������D$4��Ǆ$x     t	���0l  �3��D$Ǆ$x  �����X�L$,�QL���D$,(6�D$P�L$0Ǆ$|     �# �L$�|$���  Q��������G��~�Wi��   ��h����3�j P�L$4�# �L$��t	��Pj�ҍL$,�D$    Ǆ$x  �����S���L$$�D$P���Ec ��������L$$�4� ��u������h��V� ��2��]  �L$$�*L �\$��9��  tL��th��h��V�x h�V�m �����  ���th(�V�S h�V�H ���D$ �L$$�@ ����  �L$Q�L$(3ۉ\$��[ ;��  ��}p��t2h��V�  �D$(����=�  �D$ �>���h�V��~ ��j0�"������D$4��Ǆ$x     t	���u� �3��D$Ǆ$x  �����X�L$,�vJ���D$,(6�T$R�L$0Ǆ$|     �5! �|$�D$���  P���߹���G��~�W�@���D��3�j P�L$4�+! �L$��t	��Pj�ҍL$,�D$    Ǆ$x  �����Q���L$$�D$P���Z ��������L$$�ܭ ��u���7���hh�V��} ��2��  �L$$�RJ �\$��9��  tL��thL�h��V�} h�V�} �����  ���th��V�{} h�V�p} ���D$ �L$$�< ����  �L$Q�L$(3ۉ\$��P ;��  ��}p��t2h��V�(} �D$(����=�  �D$ �f���h�V�} ��jp�J~�����D$4��Ǆ$x     t	���M����3��D$Ǆ$x  �����X�L$,�H���D$,(6�T$R�L$0Ǆ$|     �] �|$�D$���  P��������G��~�Ok�p�D��3�3�WP�L$4�U �L$;�t	��Bj�ЍL$,�|$Ǆ$x  ������O���L$Q�L$(���|$�O ;�������L$$��� ��u���a���h0�V��{ ��2��  �\$$���zH �T$��9��  tT��th �h��V��{ h�V�{ ���D$���  �!��th��V�{ h�V�{ ���\$$�D$ ����: ����  �L$Q���D$    ��P ���  �\$ �����}e��t+hp�V�C{ �������  �����h�V�&{ ��j �l|�����D$4��Ǆ$x     t	���, �3��D$��$x  �x�L$,��F���D$,(6�T$R�L$0Ǆ$|     � �|$�D$���  P��蝷���G��~�O���D��3�j P�L$4�| �L$��t	��Bj�ЍL$,�D$    Ǆ$x  �����N���L$Q�L$(�O ��������\$ �\$$��誩 ��u�������h�V�#z ��2���  ���F �T$��9��  tP��th�h��V��y h�V��y ���D$���  ���th��V��y h�V�y ���D$ ���}9 ����  �L$Q���D$    �P ���  �
   }r��t2hX�V�sy �D$(����=�  �D$ �����h�V�Oy ��h  �z�����D$4��Ǆ$x  	   t	��腣 �3�����D$��$x  �H �L$,��D���D$,(6�T$R�L$0��$|  � �|$�D$��  P���$����G��~�Oi�  �������3�j P�L$4� �L$��t	��Bj�ЍL$,�D$    Ǆ$x  �����0L���L$Q�L$(�O ��������|$$���� ��u�������h �V�Hx ��2���  ����D �\$��9��  tL��th��h��V�x h�V�
x �����  ���th��V��w h�V��w ���D$ �L$$�$8 ����  �L$$�T$3�R�\$�xP ;��$  ��}s��t2h8�V�w �D$(����=�  �D$ �����h�V�yw ��h�   �x�����D$4��Ǆ$x     t	���/� �3��D$Ǆ$x  �����X�L$,�C���D$,(6�D$P�L$0Ǆ$|     �� �L$�|$��  Q�������G��~�Wi��   ��8����3�j P�L$4�� �L$��t	��Pj�ҍL$,�D$    Ǆ$x  �����UJ���L$$�D$P���TO ��������L$$�3� ��u�������h��V�lv ��2��  �L$$��B �\$��9��  tL��th��h��V�7v h�V�,v �����  ���thX�V�v h�V�v ���D$ �|$$���: ����  ��$�   �D$    ������$�   Ǆ$x     �a�����$�   Q�T$R���[ ����   �}?����   h�V�u �D$(����=�  �D$ ��   h�V�ju ���   �L$��(  �s1���L$,���(A���D$,(6�D$P�L$0��$|  �� �L$Q����H��j W�L$4� ��$�   R���   �p����L$��t	��Pj�ҍL$,�D$    Ƅ$x  �H����$�   �j�����$�   P�L$Q�L$,��Z ���	����L$$�#� ��u0��th��V�t ����$�   Ǆ$x  ��������2��)
  �L$$��@ �\$��9��  t-��th��h��V�Dt h�V�9t �����  �D$ ��$�   Ǆ$x  ���������"��th �V�t h�V��s ���D$ �L$$�4 ����  �L$$�T$3�R�\$�+N ;��!  ��}p��t2h��V�s �D$(����=�  �D$ �����h�V�s ��j8��t�����D$4��Ǆ$x     t	���! �3��D$Ǆ$x  �����X�L$,�&?���D$,(6�D$P�L$0Ǆ$|     �� �L$�|$��8  Q�������G��~��    +ЋG�D���3�j P�L$4�� �L$��t	��Bj�ЍL$,�D$    Ǆ$x  �����kF���L$Q�L$(���
M ��������L$$�i� ��u�������h`�V�r ��2��2  �\$$����> �T$��9��  tT��thH�h��V�Kr h�V�@r ���D$���  �!��th��V�"r h�V�r ���\$$�D$ ����3 ���k  �L$Q���D$    �XP ����   �\$ }8����   hp�V��q �������  ����h�V�q ���   �L$,�y=���D$,(6�T$R�L$0Ǆ$|     �8 �|$�D$��H  P��貵���G��~�Oi��   ��8����3�j P�L$4�+ �L$��t	��Bj�ЍL$,Ǆ$x  ������D���L$Q�L$(�xO ���$����\$ �L$$�� ��u���>���h��V��p ��2��  �L$$�Y= �\$��9��  tL��th��h��V�p h�V�p �����  ���thX�V�p h�V�wp ���D$ �L$$��4 ���  3ۍ�$�   �\$�����L$$S��$�   R�D$ PǄ$�     �Z �����@  }@����   Sh �V�
p �D$,����=�  �D$ �d���h�V��o ���   �L$$�e< �L$9��  t1��tSh��V�o h�V�o ���L$$�2< �T$���  �|$ t+�L$��X  �2,���L$��$�   �HR�H� ������+��t'��Suh�����uh��h��V�>o ����$�   Ǆ$x  ����������$�   ���D$    �M���j ��$�   P�L$ Q�L$0Ǆ$�     �zY �����������$�   Ǆ$x  �����Y����|$$���N� ��u���	���hx�V�n ��2��W  ���&; �T$��9��  tT��thd�h��V�tn h�V�in ���D$���  �!��th��V�Kn h�V�@n ���|$$�D$ ���-1 ���<  �L$Q3ۋω\$��O ����   }=����   Sh��V��m �D$,����=�  �D$ �3���h�V��m ���r���U: �T$9��  t/��tShP�V�m h�V�m �����$: �L$���  �|$ t�L$�T$R��h  ��s�����tSh�V�]m ���D$P�σ��D$    �O ���0�����脝 ���r������9 �L$��9��  tP��th��h��V�m h�V��l ���T$���  ���thx�V��l h�V��l ���D$ ���D$    �84 ����  �D$,P�L$$3�Q�ω\$(�\$4�\$8萗 ����  �|$   ��  �d/�`/�h/��$�   ��$�   �l/��$�   �D$<P�L$DQ��$�   �T$CR��$�   P�ψ\$K�\$P�\$L�1 ��ut��B���ЍL$DQ�D$(3��T$8R�ωD$<�D$L�D$P�m� ����   ��螗 ����   ��P����3�;���   w
;D$$��   �|$4  ��   3��h�L$��x  ������$�   ���$�   �P��$�   �H��$�   �P�L$@�H(�T$<�P,�L$@��P�D$@PQ���� ��t"���Q� ��t0�D$���2 ���y����/;�t+�T$Rh�V�k ���;�th��V��j ���3ۋD$�  P����� ��u���[2 ��t;�th`�V��j ���\$��S�L$P��A���L$��BǄ$x     �ЍL$LQ���n  �T$PR�K�tn  ��$�   �{�	   �t$T�{,�	   �t$x�L$L�CPǄ$x  �����ʸ �D$��$p  d�    Y_^[��$X  3��� ��]� ��R�����������U������<V��N�Lf  ��j ݞ�   ��j j ݞ�   �L$0�F    �F$   ��R��� h�   h�   h�   �L$0�F(��R���h�   h�   �N,h�   �L$0�R���0'����\$�L$@��V0�T$�$��������N8�P�V<�H�N@�P�VD�H���NH�T$�P�T$�L$@�$�VL�������NP�P�VT�H�NX�P�V\�H���N`�T$�P�T$�L$@�$�Vd�I�����Nh�P��Vl�H�Np�P�Vt�H���Nx�T$�P�T$�L$@�$�V|������$����   �P���   �H���   �P���   �H���   �Pݞ�   ���ݖ�   �L$@�艖�   ݖ�   ���T$�\$�$������艎�   �P���   �H���   �P���   �H���   �Pݞ�   ���   �F    3��F�F�F�F^��]�������������j�h�xd�    PQV�  3�P�D$d�    ��t$�S� �N�D$    �|���d  �N(�D$�M���N,�M���N0�M���N8�����NP�����Nh�������   ��������   ��������K����ƋL$d�    Y^�����������j�h�xd�    PQV�  3�P�D$d�    ��t$�|��N�D$    �Rc  ���D$������ �L$d�    Y^�����VW�|$j��j����j ����t�F P����d �����N$��  Q����d ������  ݆�   �����$�gf �����n  ݆�   �����$�If �����P  �N(Q���Cf �����:  �V,R���-f �����$  �F0P���f �����  �N8Q���1f ������   �VPR���f ������   ݆�   �����$�e ������   ݆�   �����$�e ������   ���   P����e ������   ݆�   �����$�he ����ts�NQ���c ����ta�VR���e ����tO�FP���Bg ����t=�NhQ���`e ����t+���   R���Ke ����t݆�   �����$��d ��_^� ��������̸   ����������̸   ����������̃�0SVW���L$�_����\$@S���1���wPV�D$(P����b�����P�V�H�N�P�V�H�N�P�V�w8V�D$(P���qc����L$�P�T$�H�L$�P�T$�H�L$�P�L$�T$ �������$����Au)�D$�L$�T$��D$�N�L$�V�T$ �F�N�V�whV�D$(P����b����L$�P�T$�H�L$�P�T$�H�L$�P�L$�T$ ������$����Au)�D$�L$�T$��D$�N�L$�V�T$ �F�N�V���   V�D$(P���~b����L$�P�T$�H�L$�P�T$�H�L$�P�L$�T$ ������$����Au)�D$�L$�T$��D$�N�L$�V�T$ �F�N�V_^�   [��0� �������̋A ������������̋D$�A$� �����̍A��������������D$������������z��ݙ�   � ����������{���� ����������݁�   ��$�5�$������������������D$������u��ݙ�   � ����������{���� ��V�D$����������{���$�Q�������t�D$�����ݞ�   �5ݞ�   ^� ���������̋D$�Qh��Ql�P�Qp�P�Qt�P�Qx�I|�P�H� �����̋D$���   ����   �P���   �P���   �P���   ���   �P�H� ����݁�   ���������̋D$�A,� �����̋D$�A0� �����̋I,�D$�� ���̋D$��QP�P�QT�P�QX�P�Q\�P�Q`�@�Ad� �����̋D$��Q8�P�Q<�P�Q@�P�QD�P�QH�@�AL� �����̋D$�QP��QT�P�QX�P�Q\�P�Q`�Id�P�H� �����̋D$�Q8��Q<�P�Q@�P�QD�P�QH�IL�P�H� �����̃�xV��N<�F8�V@�L$8�NH�D$4�FD�T$<�VL�L$D�L$4�D$@�T$H��������  �L$4�6�������  �L$������F$��t	����   �Nl�Fh�Vp�L$�Nx�D$�Ft�T$�V|�L$�L$�D$�T$�Q�����ta�L$�������tT�D$4P�L$��������4����Az7��$�   �L$�T$��L$�P�T$�H�L$�P�T$�H�P^��x� ������$h(��L$@�R�����t?h���D$8P�L$lQ�z�����T$�H�L$�P�T$�H�L$�P�T$ �@�D$$�=h(��L$8Q�T$lR�;�����L$�P�T$�H�L$�P�T$�H�L$ �P�T$$���L$������D$P�L$8Q�T$TR��������L$L�����L$�M����L$4�������tz�����w>�D$���D$L���������D${�D$L��P�L$�H�T$ �\$�P�L$$�T$(�p�D$�؋L$�T$�D$�D$�L$ �L$�T$$�T$�D$(�L$,�T$0�Z�D$���D$T���������D${�D$L��P�L$�H�T$ �P�L$$�T$(�\$$�H�P���T$0��A�L$,u	�L$�����L$�1���P�L$ �����������Au	�L$������$�   �L$�T$ ��L$$�P�T$(�H�L$,�P�T$0�H�P^��x� ��$�   �����������P����H����P����H�P^��x� ���������݁�   �������������D$������A{����������Az��ݙ�   � ��ݙ�   � ��������������j�hyd�    PQ�  3�P�D$d�    h�   �^�����D$���D$    t�������L$d�    Y���3��L$d�    Y������������V�t$��th�R���*����t��^�3�^����������������j�h;yd�    PQVW�  3�P�D$d�    ��h�   �a]�����D$���D$    t���������3����D$����tW���/���ƋL$d�    Y_^������������VW�|$��t5h�R����)����t%�t$��th�R����)����tW���V/��_�^�_2�^������������̋I$�����w�   � h��h��j8h���7� ��3�� ��������������̃�SUV��F$3�3ۃ�W�l$wl�$����@��   �^�,��W���   �K� ��   �?����8����   �,�   �������   �����\$������,1�|$0P�FPh��W�Z h��W�Z �NP�VT�FX�L$,�N\�L$8���L$�T$�V`�D$�FdQ�ωT$(�D$,�.] h�&W�CZ ����thp�W�1Z ���V8�N@�F<�T$�VD�L$�NL�T$ �D$�FH�T$�L$(R�ωD$(�] h�&W��Y ����thd�W��Y ���Fh�Nl�Vp�D$�Ft�L$�Nx�D$ �T$�V|�D$�L$$P�ωT$,�b] h�&W�Y ���|$ thX�W�Y �����   ���   ���   �L$���   �L$ �L$�T$���   �D$���   Q�ωT$(�D$,��\ h�&W�,Y ݆�   ��'�$hD�W�Y h4�W�Y �V(���D$0P�ωT$4�!` h�&W��X h$�W��X �N,���T$0�L$0R����_ h�&W�X h�W�X �F0���L$0Q�ωD$4��_ h�&W�X ݆�   �$h��W�zX ��_^][��� �e�e�e�e� ����+�2�^�>�L��������̃�VW�������|$�D$P�L$Q���D$    �D$    �\ �����   �|$�  �T$R���D$    �E �ȅ��Y  3�9D$�L$��Q�ωF ��D �ȅ��6  �T$R�-P �F$�����   P���YE �ȅ��  ���   Q���@E �ȅ���   �V(R���:E �ȅ���   �F,P���$E �ȅ���   �N0Q���E �ȅ���   �V8R���8E �ȅ���   �FPP���"E �ȅ���   ���   Q���D �ȅ�tq���   R���D �ȅ�t\���   P����D �ȅ�tG���   Q���zD �ȅ�t2�VR����C �ȅ�t �FP����E �ȅ�t�NQ���H �ȋT$��}B݆�   �`���������������Au���������������Au�����ݞ�   ݞ�   ��|K��t#�VhR���2D �ȅ�t���   P���D �ȃ|$|��t�Ƹ   V���C _��^��� ��_^��� ������������U����j�h�yd�    P���  SVW�  3�P��$�  d�    ��j�L$(�D$'�� �F$�����Ǆ$       ��  �$���~PW�L$(�޲����8V��$   P������P�L$(������D$,��~,�U3�9M��Q�MR�T$0QRjPj j� �� ���D$#�|$0 �t$#Ǆ$   �����D$$�$t�D$(��tj P�L$,��$�Ƌ�$�  d�    Y_^[��]� ��PV�l�����ܞ�   ������   ���ܞ�   ����A��   �~8���"����\$4݆�   ��$�5�$藾 �L$4WW��$�  �\$<�^PQ������P��$L  �n� �D$4���$P��$�  Ƅ$  �of ��$D  Ƅ$   �+ �T$TR��$�  ��f �D$$P�L$XƄ$  �& �L$TƄ$   �� ��$�  Ƅ$    �] S�o����^P��8V��$�   Q�������P�L$(����S�I�����PV�L$(�����D$# �o����~PW�L$(������hV��$`  R�����~PW�L$(�Ѱ���^hS��$�   P������P�L$(贰�����   P��$�  Q�ωD$<�j���P�L$(萰���D$4S��$0  RP��$�   Q���C������<���P�L$(�b�����$�L$4���$��$�   RS��$�   P�����������P�L$XQ���������8V��$  R�L$\�����P�L$(�	����N��V�L$@�N�D$<�F�T$D�V�L$L�L$<�D$H�T$P�7����L$4S��$H  P������������5h����L$D�$������L$<Q��$x  R�L$\������I ��a�j���a�j������������������̸�S����������������������̸�   ��������������D$������z���YP� ����������z���YP� ���\$�D$�YP� ���D$������z���YX� ����������z���YX� ���\$�D$�YX� ����V��(�77���t$%��� P���7����^� �D$�A(� �����̋A������������̋D$�A� ������V�t$��thhT��������t��^�3�^���������������̸hT�����������j�h�yd�    PQV�  3�P�D$d�    ��t$������   �D$   � �N�D$ �L  ���D$������#���L$d�    Y^����̋A$��t���t�   � �D$��th��P��O ��3�� �� �������������VW���'�����O��P  �M  _�F^��V�t$Wj j��h � @���h� ����  S�GP����O �؄���  �OQ���M �؄���  �WR���ZQ �؄��  �G!P����w �؄��i  �O$Q���M �؄��T  �W(R���jM �؄��?  �G,P���UM �؄��*  �O0Q���@M �؄��  �W4R���+M �؄��   �G8P���M �؄���   �O<Q���M �؄���   �WHR���p �؄���   ���   P���N �؄���   ���   Q���lN �؄���   ���   R���N �؄�t}���   P����q �؄�ti݇�   �����$�N �؄�tP���   Qj���qL �؄�t:��  R����M �؄�t&��   Pj���GL �؄�t��@  Q���#L �؋��
w ��u	[_��^� ��[_^� _��^� �����������̋L$3���Vw)t!��w)�$��3�ø   ø   ø   øV   Ã��u��y|�����̋L$3���wt+�t��u!�   �3�ø   Ã�t���u�ø   ��������̋L$�ɸ   t;�t
���u��3�����̋L$3���t��t���u�ø   �3��U������8SV������`/�F�d/�N�h/�V�l/3ۍN�F�^��H  �   �NH�^ �F!�F$�F(�F,�F0�^4�^8�^<�7I��j��L$@�|2���L$<���   j��L$@�g2����T$<���   �`/���   �d/���   �h/���\$���   �l/��   �$���   �F�����ݖ�   Sݖ   Sݞ�   S�  ݖ  ݞ  �V4����ݖ(  ��@  ݞ   ��ݖ8  ݞ0  �`/��D  �d/��H  �h/��L  �l/��P  ��T  ^[��]����������V�t$��thPU�������t��^�3�^���������������̸PU����������̋D$�����w7�$�(�   ø   ø   ø   ø   ø   ø   ø   �3�Ë�����������̋D$��t��t3�ø   ø   ���̋L$3�+�t��u�   �3����������j�h�yd�    PQV�  3�P�D$d�    ��t$�����  ���D$   t��Pj��ǆ�      �N�D$ �pF  ���D$���������L$d�    Y^���SU�l$��;���   ���  ��t��Pj��ǃ�      VWU����"���E�C�M�K�U�S�E�C�M�U�KR�K�M  �E �C �M$�K$�U,�S,�E(�C(�u0�{0�    󥍵�   ���   �    󥍵0  ��0  �    󥋍�  ��_^t��������  ]��[� ������SV��������  3�;�t��Pj�҉��  �`/�F�d/�N�h/�V�l/�N�F�^�/E  �N0�^ �^$�^(�E�����   �E����0  �xE���^,^[��̋Q R�w�����;�t�D$��tRh��P�H ��3�� �Q$��t��t3���   ��   ;�t�D$��t�Rh��P�MH ��3�� �I(3ҋ�+�t
��u�P�3�;�t�D$��t�QhX�P�H ��3�� �   � ������V�t$WhX�V����G ���GP���?N h�&V��G �����JG hP�V�G �G ����wW�$��hD�V�G ���Oh4�V�G ���?h �V�G ���/h�V�rG ���h �V�bG ���Ph��V�QG ��h��V�CG �O$������ t)��t��tQh��V� G ���h���h���h��V�G ��h��V��F �O(������ t��tQh��V��F ���ht��h\�V�F ��h@�V�F �����'F �O0Q����J ���UF h$�V�F ����� F ���   R����J ���+F h�V�`F ������E ��0  W���J ���F ����E _^� �c�s����������������[����  ���������D$�����D$��z	������At��������u������Au�   ��ٸ   ���������3���������U������   ��L$8�\$0�$����D$0��������0'�$����$��T$�����������2  �����������:  ��S���D$\�T$,�$P�k�����P�L$lQ��苷��� ���T$8�@�T$@�@�T$Ht6��V�؍L$<�\$,�A���� V�L$<�\$<�1����D$(��D$H�D$@�D$8������$����4���p���A�xDt,���������  ������At������At������z����������5�\$ �D$S�t$4���T$t�T$$�$R菷����P�D$TP��诶��� ���T$8�@�T$@�@�T$Ht6��V�؍L$<�\$,�e���� V�L$<�\$<�U����D$(��D$H�D$@�D$8�����%�$����4����Ata�p�������AtP�xD��������{?������At8������{3�D$ �5����DzJ���D$�M��D6��]����������������5�T$�D$ ��������Dz�M���3���]����D$���\$�$�J�������t��D$ �U��D6��]ËU����3������5���]ËU����3��5���]���̋D$��0V��P�L$Q�N0�(A���~$uV�T$<R�D$ P���   �A���D$�����D$,���������������Au�����D$���D$�D$$�����D$������D$�D$��$�L$��Q�T$ R��0  ���\$�����\$�@����L$@��P�Q�P�Q�P�Q�P�Q�@�A�~, ^�   u���Y��0� ����������U������   �EV��P�L$dQ�N0�0@���L$`藹���\$X�~$�  �UR�D$|P���   �@���D$h���L$H��Q�D$d�T$D��R�Ƀ���݄$�   ���������%�$�\$݄$�   ����݄$�   ��������݄$�   �������������\$�����������������$�� �� ��|s��t'�D$H���\$�D$P�$�!�������u�D$H�\$@�D$@�D$xP����$�   �$Q�%�����P��$�   R�L$h�@���� �T$`�@�T$h�@�\$p��D$`�D$h������������Dz��������Dz
�����T$P�����蟨 �\$P���D$p������$��D{7�ٍL$`���_����D$p���n� ��$������z���%H+���������������D$P��$�������T$`�x�������Au�������\$`�������z/�����T$`�����������������T$h������Az�����\$h�"����������z��T$`������������{����D$X�D$`P�\$t��$�   Q��0  ��=����M��P�Q�P�Q�P�Q�P�Q�@�A�   ^��]� ���U������   �ESVW��P�L$,Q�O0�~=���L$x�ů���L$(�����\$P��3��$��t$$��  �U��R�؍D$dP���   ��=����, �\$X��  �D$p��������T$X�D$8�����������������n  �������������_  �-0'�L$`Q����$�   �   �t$0�^�T$L�$R謱����P��$�   P�L$0�ǰ��� �T$x�@ݔ$�   �@ݔ$�   ����������4����At���������������������Au�����3��t$$�d$8�L$`Q���t$|��$�   �T$T�$R������P��$�   P�L$0�8���� �T$x�@ݔ$�   �@ݔ$�   ��������4����At���������������Au�����3ۅ�t)�D$H���\$�D$P�$�s�������t
�D$@�\$X��D$H���\$X�t$$����������D$0�L$H��Q�ɍT$D�D$,R�����������%�$�\$݄$�   ����݄$�   �������������\$���������$�<� �� ���h  ��t'�D$H���\$�D$P�$���������u�D$H�\$@��ua�D$@�D$`�   P�t$(����$�   �$Q輯����P��$�   R�L$0�׮��� �T$(�@�T$0�@�\$8���������������   �D$X���\$�D$P�$�9���������   �D$@�D$p���D$8�T$H�p�������A��   �xD������u|�D$h�   �ʉt$$���D$0�T$0���T$(�����������ʀ, �R  ���J  �D$8�����xD������zj�\$P����A�f  ������zD�   ���t$$��   ���؃�~�D$X�D$`P��������D$0�D$(�|����D$0�D$(�{����   �t$$�   ����� ��\$P������   �E����P�L$d��Q�؍��   ��9���D$p�����D$`����������   �D$h��������zx����������A�D$0�D$(��u�   �ʉt$$������   �ʉt$$�ɋO(���6  ��4�D$P�����ل��/  ��4�������  ��t���t�������D$0�D$(��������������������Dz��������Dz������������������+� ��������$�����5�$�T$(�x�������Au���������z�����������Au�����T$(�   9w(u���5���\$(��؀, �D$8�����T$0t4������z�����\$0�D$P��   ����������z�\$0�D$P�   �������D$P�   �D$P������Au������$�������T$(������z�����������Au�����T$(���������T$0������z�������\$0�����������Au���\$0����Ƀ�u�D$$�X+�����5�+�\$(��ٍT$(�\$8R��$�   P��0  ��6����M��P�Q�P�Q�P�Q�P�Q�@_�A��^[��]� �������������U������   �ESVW��P�L$dQ�O0�|$T�6���UR�D$|P���   �&7���L$x������   �\$X9w$�D$H    �  �, t�L$XQ�\$|�|$d�I������D$H�T$PR3��\$|�|$d�.�����9t$H��t�D$P���\$�D$h�$��������u�D$P�L$H�\$X�D$PP�   �\$|�|$d��������|$H ��t�D$P���\$�D$h�$�n�����;�u
�D$P�L$H��D$X�|$H tH�L$xQ����$�   �$R�j�����P��$�   P�L$h腩��� �|$L�T$`�@�T$h�@����   �|$L���D$`���D$h��������Az3���   �W,��t�D$p���D�`��������z�   �D�`��������Au
�L	�L$H��D	�D$H�D$x��݄$�   ��������Az3���   ��t݄$�   ���D�x��������z�   V�L$|蘬��� ������������D{������Au=�L6�L$H���D$p�D$h�D$`�������ɋt$H���H'�F�����   �$�$��������zT6�T$H���������������������F���������������8�������������*���������X+��������������������������Ƀ(��$�������T$`���������\$h�\$pu*�, t����+�������\$`�����������������؍D$`P��$�   Q��0  �^3����M��P�Q�P�Q�P�Q�P�Q�@_�A��^[��]� ��$<LZt����̋D$��0V��P�L$ Q�L$@藻���~$�T$<u7�L$HR�D$P�3���L$腬���D$@��R8P�L$Q�D$$P����^��0� �L$@�QR�P8�L$$Q����^��0� ����������̋A ���������   �$���D$P�T$R��0  �b2����L$$��P�Q�P�Q�P�Q�P�Q�@�A�   ��� �T$$�D$ R�T$ PR�������� �D$$�T$ P�D$ RP�c������ �T$$�D$ R�T$ PR�9������ 3���� �D$$�T$ P�D$ RP������� ��u9SmmmV�t$Wjj��h � @���� ��tA�GSP���x1 �؄�tW���Z3 �؄�t��W���	U �؋��@\ ��u[_^� ��[_^� �������������̃�UVWh�   3���WV�jt �N�n���E    �F�����L$�z/���D$P�L$�|$�|$�|$ Qh � @���Hj ��tz�|$S�Ä�tUU��� �؄�tGV����! �؄�t9�|$|2�t$V���  �؄�t ���K� =��}���2����t����.������] ��u
[_^]��� ��[_^]��� �V�t$Wjj��h � @���� ��tbSW���2 �؄�t?�GP���
2 �؄�t.j ���0 �؄�t�O Q����1 �؄�t�W0R����/ �؋���Z ��u[_^� ��[_^� �������������V�t$Wj j��h � @���(� ��t0SW���1 �؄�t��W����T �؋��qZ ��u[_^� ��[_^� ��������������̊A"$�����������V�t$Wj j��h � @���� ��u_^� SW����T �Ί��Z ��u2ۊ�[_^� ���������������V�t$Wjj��h � @���h� ��u_^� SW���T �؄�tL�GP����T �؄�t;�O Q����X �؄�t)�W!R����X �؄�t�G"$�D$�L$Q����X �؋��mY ��u2ۊ�[_^� ��������������̋Q2���t(�I��~!V�t$��t��~VhX  QR��� ���^� �����������̋Q2���t(�I��~!V�t$��t��~VhX  QR�u� ���^� �����������̋D$�L$i�X  PQ�[K����� �����V�t$��th�S��������t��^�3�^����������������SV�t$W���GPh�7V�8/ h`�V�-/ ���OQ���5 h�&V�/ ���O�-  ��u��7Pht7V��. h4�V��. ���W$R���6 h�&V��. h$�V��. ���G(P����5 h�&V�. hP�V�. ���O,Q����5 h�&V�. h�V�}. ���W0R���5 h�&V�d. h<�V�Y. ���G4P���{5 h�&V�@. h(�V�5. ���O8Q���W5 h�&V�. �GP��'�5��$h�V��- �GX��'���$h �V��- �GH��'���$h��V��- �G@���$h��V�- h��V�- �����   R����3 h�&V�- 3ۃ�9_l~AU3�I Sh��V�t- ������, �Gh�(�(�BV�Ћ��- ����X  ;_l|�]_^[� ���������������Q�D$��SU�ilVW�L$}3���p;�}E�\$��i�X  ��I �Ah�;X$t��u�L$��t)Q�H�+  ��t�L$����X  ;�|�_^]���[Y� _��^][Y� �������VW�|$��t5hhT���������t%�t$��thhT���������tW������_�^�_2�^�������������j�h1zd�    PQV�  3�P�D$d�    ��t$�����N�D$    ����M)  �NH�D$� %�����   ������   �������   �?�����  �D$������������ƋL$d�    Y^��������V���(����D$t	V��.������^� �̃�VW�������|$3��D$�D$�D$P�L$Qh � @��� c ���a  �|$St2��/  �VR��� �؄��  �FP���y �؄��  �NQ���T �؄���  �V!R���& �؄���  �D$P���9 �؄���  �L$Q�5������T$R�ωF$� �؄���  �D$P�_������L$Q�ωF(�� �؄��y  �T$R�y����F,���D$P���� �؄��S  �L$Q�S������T$R�ωF0� �؄��-  �D$P�M������L$Q�ωF4�{ �؄��  �T$R�'����F8���D$P���U �؄���   �L$Q�������VHR�ωF<�P �؄���   ���   P��� �؄���   ���   Q��� �؄���   ���   R��� �؄�tx���   P���� �؄�td���   Q���P �؄�tP���   Rj��� �؄�t:��  P���6 �؄�t&��   Qj��� �؄�t��@  V���l �؋���T ��u[_��^��� ��[_^��� _��^��� ������������VW�|$��t5hPU��������t%�t$��thPU��������tW������_�^�_2�^�������������j�hczd�    PQV�  3�P�D$d�    ��t$�S����N�D$    ���%  �N0�D$�@!�����   �5!����0  �*!����ǆ�      ������ƋL$d�    Y^���������V�������D$t	V�K+������^� ��SV��W�^ SjhxV4�ˁ ���;����   �F$PjW豁 �N(QjP襁 �V,RjP虁 �N0Qh�   P芁 �����  ��0��tx���t+��t��ugP��������tZ��ȋBW���LP�/ ��P�3W���؃���t7��BW���Ћˋ�������t ���   ���   P��    QW�� ������0  Vh�   W�� ��_^[�����������Vj<��j V�sh ����F4�F8���F0 ��^����������������j�h�zd�    P��SUVW�  3�P�D$,d�    ��j<3�UV�h �|$H������F4�F8�D$P�L$Qh � @���F0 �l$ �l$$�
^ ����   �|$�Ä�tV��� �؄�t�VR��� ���D$d:�l$ �l$$�l$(�ۉl$4t�D$P��� �؃|$|?��t�N Q���K �؄��V0�T$<t"�D$<P��� �؄�t�L$<Q�! ���F0���tQ ��u2�9l$(�D$4�����D$d:t�D$ ;�tUP�L$$�p:�ËL$,d�    Y_^][��$� �����������̃� �  3ĉD$S���X���L$(UVW�L$~z�@�K����D$    ~h�����    ��t$�T$�G�D$ �O��;�L$$�W�T$(�t$}&�o<�I �D$UP��<������t3����<;�|�t$�C���<;��t$|�_^]�[�L$3��a �� � �D$��t�L$VQhh�P�$ ���L$,_^][3�2��ha �� � �������̃� �  3ĉD$�D$$VP��D$�������u^�L$3��+a �� � S�^��UW~o�v�C����D$    ~]����t$�D$�O�L$ �W��;�T$$�G�D$(�t$}#�o �L$UQ��;������t3���� ;�|�t$�C��� ;��t$|�_][�^�L$3��` �� � �D$��t�T$VRh��P�# ���L$,_][^3�2��g` �� � �������V��F�V;�u>��iɘ   ��   v��|�Ky ;�}�������   ��;�}P���n���ViҘ   Vh�   j R�d �N��i��   F�����N^����j�h�zd�    P��SUVW�  3�P�D$$d�    ��t$4jj���& �؄��)  �E$P���" �؄��  �M(Q���~" �؄���   �U,R���i" �؄���   �E0P���T" �؄���   �EP�����$�*" �؄���   �EX�����$�" �؄���   j���- �؄���   j��� �؄�tj ��� �؄�tpj���� �؄�taj j j �L$$��
��P���! �؄�tDj ���` �؄�t5j ���Q �؄�t&������$�|! �؄�t������$�g! �؍L$4�  �Ml3�;ȉD$,�D$~V�}h�W$��I �:t����X  ;�|��7��|3i�X  ǋ��O�v  ��~�GP�L$8�%  3Ƀ(�����L$��t/�T$4R����" �؄�t�D$P���3 �؄�tj ���$ �؍L$4�)  ��Ul�\$3�;ЉD$~b�}h�O$�9t����X  ;�|��H��|Di�X  ǋ��O��  ��~.�GP�L$8�u$  3Ƀ(j�����L$���   �؉���\$��tF�T$4R���D" �؄�t4�D$P��� �؄�t"j ���s �؄�t�D$�����$�� �؍L$4�a  �Ul3�;ЉD$~Q�}h�O$�9Vt����X  ;�|��7��|3i�X  ǋ��O�  ��~�GP�L$8�#  3Ƀ(�����L$����   �T$4R���! �؄���   �D$P���� �؄���   j ��� �؄���   �MQ��� �؄�t{���   R���} �؄�tg�E P���,! �؄�tV�MQ���! �؄�tE�UR���J �؄�t4�E4P���� �؄�t#�M8Q���� �؄�t�E@�����$�� �؍L$4�D$,�����  �ËL$$d�    Y_^][��� �������j�h�zd�    PQ�  3�P�D$d�    hX  �������D$���D$    t�������L$d�    Y���3��L$d�    Y������������j�h{d�    PQVW�  3�P�D$d�    ��hX  �a�����D$���D$    t���������3����D$����tW���M���ƋL$d�    Y_^������������j�hK{d�    PQ�  3�P�D$d�    h�  �������D$���D$    t��������L$d�    Y���3��L$d�    Y������������j�h{{d�    PQVW�  3�P�D$d�    ��h�  �q�����D$���D$    t���g������3����D$����tW��������ƋL$d�    Y_^�����������̡`/��d/�Q�h/�A�l/V�q�Q�~ t(�F��t!�j P�B�����F    �F    �F    ^�����������̃�VW�������|$3��D$�D$�D$P�L$Qh � @����S ��t?�|$S�Ä�tV��� �؄�t��V��� �؋���G ��u	[_^��� ��[_^��� �����V��F�V;�u;������   v��|� � ;�}�������   ��;�}P���B���F��F3ɉ�H�H�H�N����F���N^����������������S�\$��U��~dW�|$��|ZV�t$��|P;�tL�E�;�B;�>�M�;�~�;�}��P����-���Ei�X  i�X  i�X  S��WV�] ��^_][� �����������QSV�t$W�����_� ��V�������_��^��[Y� j j��� �؄��  jjh � @���a� �؄���  �GP��� �؄���  �OQ��� �؄���  �WR���R �؄���  ���   P���z �؄���  �O$Q���% �؄��u  �W(R��� �؄��`  �G,P���� �؄��K  �O0Q���� �؄��6  �W4R���� �؄��!  �G8P��� �؄��  �G@�����$� �؄���   �GH�����$�x �؄���   �GP�����$�^ �؄���   �GX�����$�D �؄���   j jh � @���
� ��tp�_lUS�Ή\$�v 3�ۈD$~)3ۀ|$ t �Gh�P����� ����X  ;l$�D$|ً��,B ��]t!�|$ t�O Q���� ��t�WtR���? �G`P���JA �؄�t�OaQ���8A �؋���A ��u2�_^��[Y� ���������������j ����#+�����j�h�{d�    PQV�  3�P�D$d�    ��t$3��Fd:�F�F�F�D$�m����ƋL$d�    Y^�������������V��j ����*���D$t	V�S������^� ����������S�\$��V����   ;^��   �NW��i�X  �9�P�j �ҋFhX  �j P�=Y �N+˃���Q�SRS���%����F�Ni�X  hX  ������j R�Y �F�Ni�X  ��������R���w����F�_^[� ������������̋D$9A}	�D$��)��� ����������̋D$i�X  SUV�t$PV����2��������t,��t(;�t$W3�9{~����B���Ѓ���X  ;{|��_^][� �����������V��V2���tT�N��~MW�|$��tC��~<WhX  QR�b� 3���9~~%S3���I �F���B�Ѓ���X  ;~|�[�_^� ������������V��V2���tT�N��~MW�|$��tC��~<WhX  QR��� 3���9~~%S3���I �F���B�Ѓ���X  ;~|�[�_^� ������������VW�|$��t5h�S���
�����t%�t$��th�S���������tW���Vc��_�^�_2�^�������������SV���w���3ۉ^�`/�F�d/�N�h/�V�l/�N�F�  �N �  SSS�N$�����h�   h�   h�   �N(����SSS�N,����h�   h�   h�   �N0����h�   h�   h�   �N4�u���h�   h�   h�   �N8�^������^@S��Nd�VH�^`�VP�^a�^X�^b�^c�Y'���`/���   �d/���   �h/���   �l/���   ��t9^t�F;�t�SP�B���Љ^�^�^^[�����j�h|d�    PQVW�  3�P�D$d�    ��t$����3��N�|$�D��N  �N �D$�A  �N$�D$�����N(������N,������N0������N4������N8������~h�~l�~p�Fd0��Ft���~x�~|���   ���D$�����ƋL$d�    Y_^������������j�hI|d�    PQSVW�  3�P�D$d�    ���|$�D��wt3�9^�D$   ���t�F;�tSP������^�^�^�OdS�D$ ����%���O �D$�]  �O�\$�Q  ���D$���������L$d�    Y_^[������������������V��FW3�;�t�WP�B�Љ~�~�~_^��������������̃�V��FW3�;�t�WP�B�Љ~�L$Q�T$�~�~�|$�|$�|$Rh � @���J ��u_^��� �|$S�Ä�t
V���7 �؋���= ��u2ۊ�[_^��� �V��F�V;�u@��i�X  ��   v��|�� ;�}�������   ��;�}2P���u$���(i�X  Fj ��ȋB�ЋNi�X  NQ��������N��i�X  F���N^������j�h{|d�    PQ�  3�P�D$d�    h�   ������D$���D$    t��������L$d�    Y���3��L$d�    Y������������j�h�|d�    PQVW�  3�P�D$d�    ��h�   �A�����D$���D$    t���w������3����D$����tW���m^���ƋL$d�    Y_^������������V�������D$t	V��������^� ��SU�l$W���Ol3���~#�Wh��$;*t��t����X  ;�|������}�ٍOd�!�����|E�D$�OhV��i�X  P�L1�  �Wh�l2$�Oh�   �D1(�Wh�D20�Gh�L0Q�&����^_]��[� j�h�|d�    PQ�  3�P�D$d�    ��3�� H8�H�H�H�L$d�    Y���������������W���G�W;�uN������   v��|� @ ;�}�������   ��;�}lP����p���O����G���O_ËW���| V�t�d:t'�F��t j P���p:�F    �F    �F    �G��G��P�%\��^�O����G���O_��U����j�h}d�    P��   SVW�  3�P��$�   d�    ����u�G$�T$dP�\$p���t�  �؄��  �O(Q���_�  �؄���   �W,R���J�  �؄���   �G0P���5�  �؄���   �L$dQ����  �؄���   ���D$d������z�������������z���
���\$P�D$P�T$l�_PR�����  �؄�tu���D$l������z�������������z���
���\$P�D$P�D$O�_XP���1�  �؄�t2�L$OQ����  �؄�t �T$OR����  �؄�t�D$OP�����  �؍L$`�p�����tV�L$`Q���@�  �؄�tD�T$PR�����  �؄�t2�D$PP�����  �؄�t �L$|Q�����  �؄�t�T$|R�����  �؍L$T�=
  3��ۉ�$�   t�D$TP���$�  ��3��ۉD$X�D$\��   �L$XQ����  �؄�t}�T$\R����  �؄�tk�L$T�#
  ��u,j�L$X�D  P������i�X  Gh3Ƀ|$X�����H(�T$TR����  �؄�t �D$XP����  �؄�t�L$\Q����  �؄����\$t�'  �T$tR����  �؄��  �L$T�	  ��uJj�L$X�
  P������i�X  Gh3Ƀ|$X�������H(݄$�   �\$���   ���$�����T$TR�����  �؄���   �D$XP�����  �؄���   �L$\Q�����  �؄�t|�L$T��  ��u,jV�L$X� 
  P�������i�X  Gh3҃|$X���P(�GP����  �؄�t2���   Q����  �؄�t�W R���_�  �؄�t�GP���N�  �؃}|F��tN�OQ���g�  �؄�t=�W4R�����  �؄�t,�G8P�����  �؄�t��@W����  �����W�g!�����L$TǄ$�   �����   �Ë�$�   d�    Y_^[��]� ������SV��F3�;�t�SP�B�Љ^S�N�^�^��k����^"�^#�F �F!^[�������̃�UV��FW3�;�t�WP�B�Љ~�nW�͉~�~�k���L$Q�T$�|$�|$�|$Rh � @���F �F!�F" �F# �A ��u	_^]��� �   9D$Su9D$}2��cV���5/ �؄�tUU���� �؄�tG�|$~@�F P���? �؄�t/�F!P���. �؄�t�|$~�F"�L$$Q�ψD$ � �؋��#5 ��u2ۊ�[_^]��� ̃�SVW�������t$$3��D$�D$�D$P�L$Q���D �؄���  �D$��u�T$RV���$���_��^��[��� ����  �D$P�L$Qh � @���@ �؄���  �WR���"�  �؄��c  �GP�����  �؄��N  �OQ�����  �؄��9  ���   R�����  �؄��!  �G$P���K�  �؄��  �G(P���6�  �؄���  �O,Q���!�  �؄���  �W0R����  �؄���  �G4P�����  �؄���  U�o8U�����  �؄���  ����b =���}0������=�   u"������=�   u������=�   u�O(�M �W@R���~�  �؄��N  �GHP���i�  �؄��9  �OPQ���T�  �؄��$  �WXR���?�  �؄��  �D$ P�L$Q3�h � @�Ήl$$�l$,��> �؄���   �|$uv�T$(R�Ήl$,�d�  �؄�t�D$(P�Od�����9l$(�l$~I��$    ��t>�od�������P���� ��2����~�M��Q��������D$��;D$(�D$|����w2 ��u2��Y��tU�|$|N�W R�����  �؄�t=�|$|6�GtP���  �؄�t%�|$|�O`Q���	 �؄�t��aW���� ��]���2 ��u2�_^��[��� ������������j�hK}d�    PQSVW�  3�P�D$d�    ��t$3��H8�^�^�^�~�D$   �P;�_�_�_�F;��D$t�SP�B�Љ^S�ω^�^�5g���F �F!�^"�^#�ƋL$d�    Y_^[�����Q3���tKVPPP�D$�D$Pj j RQj �/� ��$�|$ ��th@�h4�j+h��=b ����}3�^YË�^Y�������������Q3���U�l$t���~q��tm�ɈtgW�D$�D$�D$P�D$h��  j��T$ RUVPQj 諲 ��$�|$ ��thh�h`�jJh��a ����~;�
�7 ��_]Y��. 3�_]Y�����������Q3���U�l$tf���~x��tt��~p��tl8thWf��D$�D$�D$Ph��  j��D$PUVRQj �� ����$��~;�f�~  �f�n  3��|$ th��h��j~h��a ����_]Y��̋T$SUV��L$W�m������_S�b��S��j V�wE �D$$�L$(WP������VW���0 �h���V�r����_^][� ��������V����t4��;L	t���~����uP�9�����P	�^ËP	�^ËP	�^����������V����t`��;L	tU���~�����P	�^�u��t�x ~f�  �@    ^�h$�h�h�   h���_ �P	���^ËP	�^�����������̡P	���������̋��P	������̋��t���@áL	�@����������̋�L$f�H� ��̋��t���x ��áL	�x ����̋	����t��3�9P��#ы�áL	3�9P��#ы�Ë;P	�   t��t���@�D áL	�@�D Ë���̋	����t����L	�@��~Q�L$�PQ��[ ��� �D$� �����������̋T$��t1f�: t+�	����t����L	�x ���� RQ�=� ��� ���t3Ƀ�9H����� �L	3�9H����� ��������������̋	��+P	���#�����������������VW�����t!��;L	t���~����u	P�������t$���P	�~/�L6Q�l���T6R�    �@    �p��j P��jB ��_^� ��S��V�3��t��;5L	u�D$P�q���^[� �>W�|$~AW�\������t����L	�F;�|����~Q�?Q���SVR�F ���{_^[� ;~~/�D?PV�!�����F��N��+эTR�Hj P��A ���~_^[� �������U�l$��W��~z�D$��tr�8 tmSVU�/����7�L	�ƅ�t������ޅ�t����ً@�L$P���.����C�?���ǅ�^[t�H���f�O  _]� �L	�Hf�O  _]� ��L	����t����8~�������_]� ����t���@    �_f�  ]� ���@    �_f�  ]� ���SVW�|$����~e�\$��t]f�; tWW�O�����?PSQ�D ��L	����t������x�6�ƅ�t�P���_f�V  ^[� ���P_f�V  ^[� ��L	����t����8t�������_^[� ����t���@    �_^f�   [� ���@    �_^f�   [� ����SU�l$�����   �D$����   �8 ��   ���t����L	�@VW�P�^�����L	����t���������t�����Ѕ�t����ыȅ�t����L	�R+Q�v�L$R�4p���6���G�������_^t���@]f�A  [� �L	�@f�A  ][� ��VW�|$������   S�\$����   f�; t|���t����L	�@U�P������-L	����t����ŋ@�?R�ASQ��B �����t�����x�6�ƅ�t�P�]��[_f�V  ^� �ŋPf�V  ][_^� ����������̋T$�ҡP	V��t#�: t��W�x�I �����u�+�RP������_��^� ����̋T$�ҡP	V��t'f�: t!��W�x��f���f��u�+���RP���8���_��^� ̡P	VW�|$����~AW����3���~f�L$�f�B��;�|�f�x  ���t���x_��^� �L	�x_��^� �����U�l$V��M 9�  �L	����t����x ���-����P	���^]� ����t����8 ~C�8 ��u4��������E ��t��� �M ���^]� �L	� �M ���^]� �L	�E ��t����PSR�������M �L	����t����Ëх�W�xt�����3�9B�?��R��#ȋQP�@ �E ����_t����Ë�ɋ@t��[�A��^]� �ˉA[��^]� ��������̋T$W��;t,��t��V�p�����u�+ƍH������^v3�RP��������_� ��̋T$W��;t0��t!��V�pf���f��u�+����H������^v3�RP���%�����_� ���������������V�D$Pj��������^� �����������V�t$��W��t�ƍP�����u�+H������v3�VP��������_^� �������V�t$��W��t�ƍPf���f��u�+����H������v3�VP��������_^� ��́�  �  3ĉ�$   VW��$  h   �D$j P�; ��$   ����t#��$  QP�T$h�  R�l� ��Ƅ$   �D$�P�����u�+��F�=���w��}&���w����P	�_^��$   3���5 ��  �V���0����T$RV���������$  _^3���5 ��  ������������̸  ��B �  3ĉ�$   VW��$  h   �D$j P�.: ��$   ����t%��$  QP�T$h�  R�� ��fǄ$    �D$�P�d$ f���f��u�+������F�=���w��}&�������P	�_^��$   3��5 ��  �V���B����T$RV���������$  _^3���4 ��  ���������������SVW������tM��;5L	tB��t>�>~9�
����P	��NSQ���g����F;F}�?��t
���G_^[Ë=L	�G_^[���V�t$���W��t����L	�8 ~/��� ��u&�����t��� ��_^� �L	� ��_^� �P	��6;�t.��t�ƍPf���f��u�+����H������v3�VP��������_^� ��W���L$����;t2��t#��V�q��    �����u�+΍Q������^v3�PQ��������_� ��������V����Wt����L	�|$;x|W������|E���t����L	;x0���}������t���x�f�x  _^� �L	�x�f�x  _^� ���������������V���8����6�ƅ�t��3�9H����#΋�^áL	3�9H����#΋�^�������SW����Å�t����L	�x �%  �|$ u�D$\��U3�f���  �D$V�0f���L$t��f;�t�A��f��u��f�9 t�����if��uͅ���   f�<k ��   ���tJ��;5L	t?��t;�>~6�������P	��FSP��������N;N}���t����L	�H��i�f�����f��u���t^��)h]_[� �L	)h^]_[� �Å�t!��;L	t���~����u	P�X�����P	�^]_[� ������QU�)�Ņ�V�L$t����L	�p����   S�\$��u�\���Wx2�|u �d$ �f��t�f����tR��f;�tJ�A��f��u��}L�Ņ�t!��;L	t���~����u	P������P	�L$_[^�]Y� f�9 t�������}��f�|u t8�L$������D$�f�Dr  � ��t_����[�p^]Y� �L	���p_[^]Y� ��VW�|$W�������W������_^� �����V�t$��th@V��������t��^�3�^���������������̸@V������������5�����D{4�Q����D{*�Y����D{"�j���%�$����'����Az�   ���3�����������A�H�����A�H������'����Az�   �3�������x���SV��ݞ  3��x��D$ݞ   P��(��V�F�^ �F	��'�^
�^(�^�F   �^�^�^�^��g����N0�P�V4�H�N8�P�V<�H�N@�P�VD���FH���NL���VP���FT� ��NX�$��V\����F`����Nd� ��Vh���Fl���Np���Vt���Fx���N|�����   �����   � ����   �$����   �(����   �,����   �0����   �4�������   �8����   �<�ݖ�   �����  ݖ�   ��  ݞ�   ���   ���   ݞ�   ���   ݆  ���   ݞ�   ���   �p����   ݞ�   ǆ�      �������  �~���������   ������   ������   ������   �����   �����  �`/��  �d/��  �h/��  �l/��  ^[�������j�hx}d�    PQV�  3�P�D$d�    ��t$� �N�D$    ����`���N0�`���NH�}`���N`�u`���Nx�m`�����   �b`�����   �W`����  �������  ������������ƋL$d�    Y^��������������u �����SU�l$��;���  VWU�x����E�C�M	�K	�U
�S
�E�C�M�K�U�S�E�C�M�K�U�S�E�C�M �K �U$�S$�E(�C(�M,�K,�U0�S0�E4�C4�M8�K8�U<�S<�E@�C@�MD�KD�UH�SH�EL�CL�MP�KP�UT�ST�EX�CX�M\�K\�U`�S`�Ed�Cd�Mh�Kh�Ul�Sl�Ep�Cp�Mt�Kt�Ux�Sx�E|�C|���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ݅�   ݛ�   ��  ݅�   ��  ݛ�   ݅�   ݛ�   ݅�   ݛ�   ݅�   ݛ�   ݅�   ݛ�   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ��   ��   ��  ��  �    󥍵�  ���  �    �݅   ݛ   ݅  ݛ  ��  ��  ��  �H��  �P��  �@_��  ^]��[� ̀y u�D$��thP�P�� ��3�� �y	 u�D$��t�h,�P�� ��3�� �y
 u�D$��t�h �P�u� ��3�� �   � ����̃�0W���	 ��   � ��   ݇�   SV���   V���D$�$P��U_����P�L$(Q�O�^����L$@��P�Q�P�Q�P�Q�P�Q�@�A�W`�Q�Gd�A�Wh�Q �Gl�A$�Wp�Q(�Gt�A,�Wx�Q0�W|�Q4���   �Gx�Q8�P�Q<�P�Q@�@�AD��QH�F�AL�V�QP�F�AT�V�QX�F�A\�(/ ^��[_��0� 2�_��0� ���̃�0W���	 ��   � ��   ݇�   SV���   V���D$�$P��U^����P�L$(Q�O�]����L$@��P�Q�P�Q�P�Q�P�Q�@�A�W`�Q�Gd�A�Wh�Q �Gl�A$�Wp�Q(�Gt�A,�Wx�Q0�W|�Q4���   �Gx�Q8�P�Q<�P�Q@�@�AD��QH�F�AL�V�QP�F�AT�V�QX�F�A\�(. ^��[_��0� 2�_��0� ����VW��� t�w���d����t�L$V�`��_^� �t$h�����	]����t���~d����u_^� ��G�V�O�Q�F�A�V�Q�F�A�V�Q�Jd����u�G�G_^� ����������́�   SV��^0W���F �d�����  �~H���d�����  �L$<�$Z���L$�Z���L$$�Z���~ ��   �~ ��   �O��W�L$�O�D$�G�T$�W�L$�L$�D$�T$ �c������   �L$�a������   �D$P����[���L$Q����$�   �$R�/\����P�D$pP�L$\Q���z^�����C[����T$$�H�L$(�P�T$,�H�L$0�P�T$4�@�L$$�D$8�c����t�L$$�`������   _^2�[�Đ   ÍL$TQ���^����T$$�H�L$(�P�T$,�H�L$0�P�T$4�@�L$$�D$8�b����t��L$$�5`����t��L$$Q����Z���T$$R���D$`�$P�P[����P�L$pQ���Z����T$�H�L$�P�T$�H�L$�P�T$�@�L$�D$ �>b�����:����L$�_�����)����L$$Q�T$R�D$\P��a����L$H�P�T$L�H�L$P�P�T$T�H�L$X�P���L$<�T$P��a����������L$<�[_����������L$<�*�����������L$������������L$$������������D$�L$<�C����������D$$�L$�.������j����D$<�L$$�������U����D$<�L$@�T$D�F`�D$H�Nd�L$L�Vh�T$P�Fl�D$�Np�L$�Fx�D$�N|�L$�Vt�T$���   �T$ ���   �D$$���   �L$(���   �D$0���   �L$4���   �T$,���   �T$8���   ���   �N���   �`��_�F^[�Đ   ËD$�Q��Q�P�Q �P�Q$�P�Q(�I,�P�H� �����̋D$�Q0��Q4�P�Q8�P�Q<�P�Q@�ID�P�H� �����̀|$ t�I� �a�� ����������̀|$ t�I� �a�� ����������̋D$��t�A��A �X�A(�X�D$��t�A`��Ah�X�Ap�X�D$��t�Ax�݁�   �X݁�   �X�D$��t݁�   �݁�   �X݁�   �X�A� ������̋D$�Q`��Qd�P�Qh�P�Ql�P�Qp�It�P�H� �����̋D$�Qx��Q|�P���   �P���   �P���   ���   �P�H� ���������̋D$���   ����   �P���   �P���   �P���   ���   �P�H� ���̋D$;Au�� ��u��A   � �����A   � ̋A�������������3��y��������̃yu�y t�I��t��u��2����D$SV���$��2��M��������  �D$���$��L��������  �D$$���$��L��������  �D$���$�L��������  �D$,���$�L��������  �D$4���$�L�������l  �D$�D$�������S  �D$$�D$�������&  �D$,��$����A�  �D$4������A�  �~ul��&������t���@�������zL��h����h����h�  ��h�������? �D$���D$�D$�D$4�D$$�D$,�����������ʊN��$��t%����������D{��������������������������tR����������D{E�������������������F	ݞ�   ���ݞ�   ݞ�   ݞ�   ��ݞ�   ݞ�   ^[�0 ������������������
������������ht�h��h�  h����> ��^��[�0 ��������������̋D$��t݁�   ��D$��t݁�   ��D$��t݁�   ��D$��t݁�   ��D$��t݁�   ��D$��t݁�   ��A	� ���������̋D$��t���   ��D$��t���   ��D$��t���   ��D$��t���   ��D$��t���   ��D$��t���   ��A
� ���������̃�V���   +��   ���   +��   �~
 �D$�D$�L$�\$�D$�T$tE���$�I������t5�D$���$�I������t�����D$��������D{�|$������������T$��~
 ^t������D{�   ��� ����3���� �����������̋T$��0��t=��D$(P��D$P�D$(P�D$$P�D$ P�D$P�.�����t���$������Az����2���0� �D$���D$������Au������D$���D$ ������Au�����������t�p�����u�������������A{��h�������0� ���������U�����E��<V���$���fH��������   ���]������   �D$8P�L$Q�T$8R�D$4P�L$0Q�T$,R���F�����tz���D$��������A{g�D$�����D$ ������Au��������D$(�����D$0������Au�������������t������u�������������u������������2�^��]� ���u�h��������%�$����'����z�ڰ����������^��]� ��0�͋������������D$h�\$(���\$ �\$���\$���\$�$����^��]� ������S�\$��UVW��t��l$��t�] ����  ���$���*�������   ݆x  ����������D��   ݆�  ������D��   ݆�  ������D��   ݆�  ��$����D��   �݆@  ��;������z_������zX݆   ������DzI݆(  ������Dz:݆8  ������Dz+݆H  ��������Dz'��t���؅�t_�] ^][� ��_��^��]��[� ����_^][� ��������������V��L$�$W����u�D$P����R����u^� �L$�T$���   �L$���   �T$���   �L$���   �T$��   ��  �^� ������̋D$���   ����   �P���   �P���   �P��   ��  �P�H� ����U������4�5SV�T$��~ W��   �]�؄�t�~	 u2ۍ��   ���@V����tU���   PW�L$0Q�N�WN�����N���T$ ����   ���$��D������t���D$ ��������Az���5��D$ ��t~���5��������Dzi݆�   ܞ�   ����AzV��݆�   ܆�   ��$ܖ�   ����z
��݆�   �ܖ�   ����Au��݆�   ��������t��_^[��]� ��_^[��]� ��������j�h�}d�    PQ�  3�P�D$d�    h(  �������D$���D$    t���k����L$d�    Y���3��L$d�    Y������������j�h�}d�    PQVW�  3�P�D$d�    ��h(  �������D$���D$    t����������3����D$����tW�������ƋL$d�    Y_^������������VW�|$��t5h@V���*�����t%�t$��th@V��������tW���F���_�^�_2�^�������������V������� �D$t	V���������^� ������������U������4SVW�������}�D$8P�L$@Q���D$D    �D$@   �i�  �؄��  �|$<�t  �T$4R���D$8    �`�  �؄���  �|$4 �L$4��Q�ψF�?�  �؄���  �|$4 �D$4��P�ψV	��  �؄���  �|$4 �T$4���N
R�����  �؄���  �D$4P�y� ���NQ�ωF��  �؄��v  �V0R����  �؄��a  �FHP����  �؄��L  �N`Q���y�  �؄��7  �VxR���d�  �؄��"  ���   P���L�  �؄��
  ���   Q�����  �؄���  ���   R�����  �؄���  ���   P����  �؄���  ���   Q����  �؄���  ���   R����  �؄���  ���   P���l�  �؄��z  ���   Q�����  �؄��b  ���   R����  �؄��J  ���   P����  �؄��2  ���   Q���|�  �؄��  ���   R���d�  �؄��  ���   P���L�  �؄���   �|$8��   ��  Q���I�  �؄���   �|$8��   �T$0R���D$4 �c�  �؄�t�|$0 ���F���D$0 t�L$0Q���=�  �؄�t�|$0 �V���D$0 t�D$0P����  �؄�t�|$0 ���N���D$0 t�T$0R�����  �؄�t�D$0P���_������D$0 t�L$0Q�����  �؄�t�T$0R���X����~ tD�N�jP����t�NH�^P����t�N0�RP����u h��h��h�  h����2 ���F �~	 �  ݆�   ���$��>��������   ݆�   ���$�>��������   ݆�   ���$�>��������   ݆�   ���$�>������tx݆�   ���$�g>������t`݆�   ���$�O>������tH݆�   ܞ�   ����t5݆�   ܞ�   ����t"��ܞ�   ����t݆�   ܞ�   ����u hP�h��h�  h���1 ���F	 _^��[��]� ����U������4SVW�}j��j����  ����  3�8F����P��  ��3�8F	����t
P����  ��3�8F
����t
P����  �؋F�ωD$<��� ��
�   9Ft�D$<����  P���]�  �؄���  �NQ���(�  �؄���  �V0R����  �؄���  �FHP�����  �؄��x  �N`Q�����  �؄��c  �VxR�����  �؄��N  ���   P����  �؄��6  ݆�   �����$�_�  �؄��  ݆�   �����$�B�  �؄���   ݆�   �����$�%�  �؄���   ݆�   �����$��  �؄���   ݆�   �����$���  �؄���   ݆�   �����$���  �؄���   ���   Q����  �؄�tt���   R����  �؄�t`���   P�����  �؄�tL���   Q�����  �؄�t8���   R�����  �؄�t$���   P����  �؄�t��  Q����  �؄ۊV�T$<t�D$<P�����  �؄ۊN�L$<t�T$<R����  �؄ۊF�D$<t�L$<Q����  �؊V����ۈT$<t�D$<P���u�  �؊N���ۈL$<t�T$<R���Y�  ��_^[��]� _^��[��]� �U����j�h~d�    P���   SV�  3�P��$�   d�    ��L$D� �D$DP��Ǆ$      �����؄��m  ��L$$Q�T$ �T$ �\$(R���H������D$�����D$<�L$T�T$,���t$4�T$4܎�   �\$܎�   �$P� ��M��P�Q�P�Q�P�Q�P�Q�@�A݆�   �L$$���L$<�\$݆�   �L$,�$Q�L$X�� ��M��P�Q�P�Q�P�Q�P�Q�@�A݆�   �L$$���L$<�\$݆�   �L$,�$Q�L$X�| ��M��P�Q�P�Q�P�Q�P�Q�@�A݆�   �L$$���L$<�\$݆�   �L$,�$Q�L$X�+ ��M��P�Q�P�Q�P�Q�P�Q�@�A�L$DǄ$   ������ �Ë�$�   d�    Y^[��]� ���������U����j�h;~d�    P���   SV�  3�P��$�   d�    ��L$D� �D$DP��Ǆ$      �����؄���  �~��u݆�   ܶ�   �\$$��T$$�L$�T$Q�\$�T$ R���,������D$�����D$<�L$T���t$$�D$4�����T$$�����T$,݆�   �����\$܎�   �$P�� ��M��P�Q�P�Q�P�Q�P�Q�@�A݆�   �L$���L$<�\$݆�   �L$,�$Q�L$X� �D$��M��P�Q�P�Q�P�Q�P�Q�@�A܎�   ���L$<�\$�D$,܎�   �$Q�L$X�P ��M�D$��P�Q�P�Q�P�Q�P�Q�@�A܎�   ���L$<�\$݆�   �L$,�$Q�L$X�� ��M��P�Q�P�Q�P�Q�P�Q�@�A�L$DǄ$   ������ �Ë�$�   d�    Y^[��]� ������������́��   SVW��|$�   ���>������y�D$TP�L$@Q�T$,R�D$P��������t$��$�   Q��$�   R��$�   P�L$xQ���j������V�N��$�   �V ��$�   �N$_��$�   �V(��$�   �N,^��$�   ��$�   [t2��$�   ��$�   3�9�$�   ��RPQ�T$Rjj	j j�Ȓ �� �����   � ���������V��~ Wt4�~0����F����t&��;�����$�E����u�L$W�GB��_^� �|$���F����tF��;�����$�`E����u/��F0�O�N4�W�V8�G�F<�O�N@�W�ΉVD�B���_^� _2�^� ������V��~ Wt4�~H���LF����t&��;�����$��D����u�L$W�A��_^� �|$���F����tF��;�����$��D����u/��FH�O�NL�W�VP�G�FT�O�NX�W�ΉV\����_^� _2�^� ������U�����E��t  S�]@;CVWt3Ƀ������K�E8�p����M<|��|	�E<�\$(��T$(��|
��|���E8��$�  �\$0�������$   �������$   �������$�   ��������T$(����Au��2�_^[��]��\$0����At����U(����t��]0����t֋�=�E��=���ĉ� >�H�>�P�>�H�>�P�(��H�,����ĉ�0��H�4��P�8��H�<��P�H����$�  �$������E��=��=���ĉ� >�H�>�P�>�H�>�P����H������ĉ� ��H���P���H���P�H����$8  �$�7�����=��=���ĉ� >�H�>�P�>�H�>�P�H���(��E �,��ĉ�0��H�4��P�8��H�<��P�H����$8  �$������$�  R��$�  P��$  Q��$  R��$  �"�����������    ��$�   h��D$<�P��$�   ����P�������L$8Qh(��T$XR��$�   �r������>��P��������D$PP���W����E0P���L$D�$Q�;���u��P�T$lR����:��P���������V���ĉ�P�N�V�H�N�P�V�H�ˉP�:����E0�������������z��������H'�D$(�D$0�����E(��A��z�������������{u�������˃�0���\$(�����\$ �T$���\$�T$���$�����D$(�� �D$0���� 3�;�t0;�t,���   ���   ���   ���   ���   ǃ�   ��  �C
��PQ����_��^��[��]������������U������8V�uWh�V���� �����{� h �V��� �G����t��th���h���h��V��� ��� �tEu�lEPh��V�� ������ h�LV�� ��� th��V�� ���GP���Q� h�&V�f� h��V�[� ��� th��V�G� ���O0Q����� h�&V�.� h(gV�#� ��� th��V�� ���WHR����� h�&V��� h��V��� ���G`P���� h�&V��� h��V��� ���OxQ���y� h�&V�� h��V�� �����   R���R� h�&V�� �����=� h��V�r� �����   P���A� h�&V�V� ��j���*������$hp�V�9� ��O	�T$H����t+݇�   ܧ�   ��������D{݇�   ܧ�   ���\$8��؄ɸtEu�lEPhL�V��� �����X� �G�tEu�lEPh(�V�� ���G�tEu�lEPh�V�� h��V�� ݇�   �����$�� h�&V�t� h��V�i� ݇�   �����$�� h�&V�K� h��V�@� ݇�   �����$�m� h�&V�"� h��V�� ݇�   �����$�D� h�&V��� h��V��� ݇�   �����$�� h�&V��� h��V��� ݇�   �����$��� h�&V�� h��V�� �D$H�����$��� h�&V�� ���u\����� ݇�   ܷ�   ���$h��V�S� ݇  ���$h��V�<� ݇   ���$hd�V�%� ������� ����� ��L$8�\$8Q���"����
 �tEu�lEPhH�V��� �����\� ���   Rh<�V��� ���   Ph0�V�� ���   Qh$�V�� ���   Rh�V�� ���   Ph�V�� ���   Qh �V�p� ��Hh��V�b� �D$@���$�� h�&V�I� ������� ����� _^��]� ��  V���F����  �F�N�V S�D$8�F$U�L$@�N(�D$H�FHW�T$H�V,�L$PP��$�   �T$X�D$`�J3���F0P��$�   �D$d�63���F`P��$  �D$\�"3���^xS��$�   �3�����   U��$�   ��2����$(  �D$@P�L$hQ��跿���T$dR�D$,P��$�   Q��$�   R�L$P�3��P��$�   P��脿������3���L$dQ�T$R��$�   P��$�   Q�L$P�z3��P��$�   R���J������3���~ t*�F�N�V �D$d�F$�L$h�N(�T$l�V,�D$p�L$t�T$x�~ t)��K�S�D$(�C�L$,�K�T$0�S�D$4�L$8�T$<�~ t5�D$|P���"6����L$�P�T$�H�L$�P�T$�H�L$ �P�T$$�L$(��:�����  �L$�:�����  ��;���L$0�$�R9������  ��;���L$�$�59������  ��;���$�D$P�L$4Q��$�   R�
:������� 9������  �F��tg�~ ug�L$�7���D$(P�L$�t2������;����A��   �L$|Q���%5����T$�H�L$�P�T$�H�L$�P�T$ �@�D$$�Y�~ tS��uO�L$(�G7���L$(Q�L$�	2������;����Az)��C�K�T$(�S�D$,�C�L$0�K�T$4�D$8�L$<�~ u�T$dR�������~ u�D$P���M����~ u�L$(Q�����������������u{�T$@�D$D�L$H�V�T$L�F�D$P�N �L$T�V$�F(��$�   �N,�L$\R�0���L$`��$�   P��/����$  Q�L$\��/����$�   R����/����$�   P����/����_][^��  � _][3�^��  � ������V���^�N�   �J�����^�������VW�|$W���b� �����tPj谮 �^���N�2���_��^� ����������̃������������̃���UV��N�^�nW�   �L$�����|$ 3��D$�D$�D$P�L$Qh � @���*�  ��u	_^]��� �|$�S�ÄۉT$t=�D$P��莪  �؄�t+�L$Q螬 ��U�ω��  �؄�t�T$R���O�  �؋����  ��u2ۊ�[_^]��� ����V�t$Wj j��h � @���\ ��u_^� �SP����  �؄�t#�G�����$螼  �؄�t��W��蝾  �؋����  ��u2ۊ�[_^� ������j�hh~d�    PQVW�  3�P�D$d�    ��L$蒹������D$    �L  �$�`�h���@  h���6  h���,  h���"  h���  h���  h���  h����   h����   h����   hx���   hl���   h`���   hT��   h<��   h4��   h,��   h$��   h��   h��   h���{h���th���mh���fh���_�~��蓸����~/���ظ����tOf�8 tI�F���$P�D$h��P�u������+�F���$�L$h��Q�X������ht��L$�����L$�������t�T$ Ph`�R�غ ���L$�D$���������L$d�    Y_^��� Ȓ����,�J�T�^�h�|���Ғܒ���"�6�@�r���������������������Vj��薩 Pj��� �^���N�N�����'�^�F0    �P<�F4   �^ ���p&�^(^��SV�t$W��jf����  �؄ۋtLP����  �؄�t>�G�����$蘹  �؄�t(�G �����$肹  �؄�t�G(�����$�l�  �؄ۋG0t
P��軷  �؋G4��|��~!h8�h�hh  h���D ���   ��t1P��耷  ��t'�G�����$��  ��t��W����  _^[� ��_^[� ������������������SV��3�S3���F   �FX  �^f�FS�F�^S�N�F   �C���h�   h�   h�   �N$�^ �)���h�   h�   h�   �Nh�����N(�ڴ���@'�   �^`�^,�^0�^4�^<�^@�^D�^H�^L��  �^n�^o�^r�F8�FP�FT�NX�N\�Fl�Fm�Fp�Fq�Fs�Ftf�^u�^w^[������������j�h�~d�    PQV�  3�P�D$d�    ��t$�N�����N$�����N(�����Nh�D$    �Н����������ƋL$d�    Y^���������j�h�~d�    PQV�  3�P�D$d�    �L$�q(���D$    �ȳ�����D$����蹳���L$d�    Y^�����������SV�t$W��jg���~�  �؄���   �P���j�  �؄���   �OQ���U�  �؄���   �WR���@�  �؄�ts�GP���߶  �؄�tb�O Q����  �؄�tQ�W$R��轶  �؄�t@�G(P��謸  �؄�t/�O,Q����  �؄�t�W0R���ڴ  �؄�t�G4P���ɴ  �؋�� ~ ��|�G8��   ����   P��衴  �؄���   �O<Q��茴  �؄���   �W@R���w�  �؄���   �GDP���b�  �؄���   �OHQ���M�  �؄�t}�WLR���<�  �؄�tl�GPP���+�  �؄�t[�OTQ����  �؄�tJ�WXR���	�  �؄�t9�G\P�����  �؄�t(�G`�����$肵  �؄�t�G�����$�l�  �؄ۋGt-P��軳  ��t#�OhQ���\�  ��t�WR�����  _^[� ��_^[� ��������������QSVW���5����|$�D$P���D$    �]�  �؄��$  �L$�����c�  V���;�  �؄��  �VR���&�  �؄���  �FP����  �؄���  �NQ��蜢  �؄���  �V R����  �؄���  �F$P���r�  �؄���  �N(Q��警  �؄���  �V,R��訡  �؄��o  �F0P��蓡  �؄��Z  �N4Q���~�  �؄��E  �V8R���i�  �؄��0  �F<P���T�  �؄��  �N@Q���?�  �؄��  �VDR���*�  �؄���   �FHP����  �؄���   �NLQ��� �  �؄���   �VPR����  �؄���   �FTP���֠  �؄���   �NXQ�����  �؄���   �V\R��謠  �؄�tw�F`P���+�  �؄�tf�|$e|_�NQ����  �؄�tN�T$R���q�  �؄�t<�D$P聢 ���|$f�F|%�NhQ����  �؄�t�|$g|��V��葮  ��_^��[Y� �����̃�d�(�����������VWjh3���WV�Q� ������V�Nd�V�~H�V�~L�V �~P�V(�~T�^0�~X�~\�~`�ۮ�����V8_�^<�F@�FA^��������̃�SVW�������|$ �D$P�L$3�Q�ω\$�\$�d�  �|$��  9\$��  ���  V����  ����   �VR���ܟ  ����   �FP���ɟ  ����   �NQ��趟  ����   �V R��裟  ����   �F(P��萟  ����   �N0Q���}�  ����   �T$ R���ٞ  ��tu�D$ P�� ���NLQ�ωFH躞  ��tV�VPR��諞  ��tG�FTP��蜞  ��t8�NXQ��荞  ��t)�V\R���~�  ��t�F`P���o�  ��t�NdQ���P�  �|$U�n@�] �^A� ��   ���F8�\$tF�T$R�����  ��t6�D$���$��������t���D$��������u�^8���U���7�  �|$|a���F<�\$tV�D$P���i�  ��tF�D$���$�������t(���D$��������uS�^<����  ]_^[��� ��S���ϛ  ]_^[��� _^2�[��� ����������U������4SV�uWj��j����  �؄���   ������$�ۯ  �؄���   �G�����$���  �؄�tj�G�����$諯  �؄�tT�G�����$蕯  �؄�t>�G �����$��  �؄�t(�G(�����$�i�  �؄�t�G0�����$�S�  �؄ۋGHtNP��袭  �؄�t@�GLP��葭  �؄�t/�OPQ��耭  �؄�t�WTR���o�  �؄�t�GXP���^�  �؋O\�L$<���v ��)�G\��t��t
�D$<    ��D$<   ��D$<   ��t0�T$<R����  �؄�t�G`P�����  �؄�t�OdQ��螰  �؄��G8t#�����$�x�  �؄�t�W@R��薪  ����؄��G<t&�����$�L�  ��t�GAP���l�  _^[��]� �؊�_^[��]� ������j�h�~d�    PQV�  3�P�D$d�    ��t$���   �D$    �U������D$�����&f �L$d�    Y^��������SV��W���   � �������    �hY�ݓ�   ݛ�   _^ǃ�   F   ǃ�      ƃ�   [������VW�|$j��j���}�  ��tV����  ��ts݆�   �����$�:�  ��t\݆�   �����$�#�  ��tE���   P���q�  ��t3���   Q���_�  ��t!���   R�����  ��t���   P���z�  _^� ����̃�SU��V���   W�L$ �(����荅�   �D$�    �hY���ݕ�   ݝ�   �t$,� F   ���   �D$�    ���   �D$$� 3��D$�D$�D$P�L$���   Q���   ��脰  ��tn�|$ugU���њ  ��tDW����  ��t8S���	�  ��t,�T$R���i�  ��t�D$P���Y�  ��t�L$ Q���9�  �|$|��t�T$$R��蒧  _^][��� ��������VW�|$j ��j���ͯ  ��tn������$蚫  ��t[�F�����$膫  ��tG�FP���ש  ��t8�NQ���ȩ  ��t)�VR��蹩  ��t�FP��誩  ��t�N Q��蛩  _^� �����̃�VW�|$��D$P�L$Q���D$    �D$    �D�  ��ti�|$ubV����  ��tV�VR���Ҙ  ��tG�FP���3�  ��t8�NQ���$�  ��t)�VR����  ��t�FP����  ��t�� V�����  _^��� ���������������SV�t$W�����r 3ۃ��Ë�Sj�~�  ��to�G P��诨  ��tK������$�<�  ��t8�G�����$�(�  ��t$�G�����$��  ��t�G�����$� �  ��|��t�O$Q����  _^[� �����U������SV3�W�}�D$�D$��D$P�L$Q�����  ����^��V��Ȅ�����F�ɉT$��D$�F     �F$ �F% �F& �F' tx�|$uq�F ��P�؋����  �Ȅ�tTV���B�  �Ȅ�tFS���4�  �Ȅ�t8�T$R���"�  �Ȅ�t&�D$P����  �Ȅ�t�|$|�F$P��訔  ����T$��������z�����������Au��������Az�������Az�������t$������z�����������Au��������Az���������Az����_^[��]� _��^��[��]� ����j�h(d�    PQV�  3�P�D$d�    ��t$���   �D$    蕤�����D$�����f` �L$d�    Y^��������VW�|$j��j����  ����   ���   P����  ��to݆�   �����$���  ��tX݆�   �����$詧  ��tAV�����  ��t5���   Q���*�  ��t"���   R����  ��t���   P����  _^� ��������������̃�VW�|$��D$P�L$Q���D$    �D$    �d�  ����   �|$��   ���   R���S�  ��t,���   P����  ��t���   Q���ϔ  ��tV���s�  �|$|N��t���   R���z�  �|$|5��t���   P���a�  �|$|��t�Ɩ   V���H�  _^��� 2�_^��� ������VW�|$j��j���}�  ��t(V���a�  ��t�FP�����  ��t�NQ�����  _^� �����������̃�SUVW��肢���|$3��D$�D$�D$P�L$Q�n�^���E � �&�  ��t8�|$u1V���#�  ��tU��臡  �|$|��tS���t�  _^][��� 2�_^][��� �������������̃�8�������������V�t$Wj j��h � @���HE ��u_^� �SP��责  �؄���   �G�����$�:�  �؄�t{�G�����$�$�  �؄�te�G�����$��  �؄�tO�G �����$���  �؄�t9�G(�����$��  �؄�t#�G0�����$�̤  �؄�t��8W���˦  �؋���  ��u2ۊ�[_^� ���̃�V�t$3�W�D$�D$���D$P�L$Qh � @���E�  ��u_^��� �|$S�Ä���   W��谑  �؄�ts�WR���/�  �؄�tb�GP����  �؄�tQ�OQ����  �؄�t@�W R�����  �؄�t/�G(P����  �؄�t�O0Q���ڑ  �؄�t��8W���)�  �؋���  ��u2ۊ�[_^��� ��������������̃�0SUV��W��X  �����������D$P���I������@  �P��D  �H��H  �P��L  �H��P  �P���  ���   ��T  賟����    �hY���ݓ�   ݓ�   ��ǃ�   F   ǃ�      ƃ�   �`/��\  �d/��`  �h/��d  �l/��h  ǅl     3����  ��ݕp  ���  ݝ�  ���  ���  ݕx  ���  ݝ�  ���  �m�����u"�L$Q��謽��P�T$,R���o���PS���� ��  ƅ�  ƅ�  ƅ�  �    �hY���ݓ�   ݛ�   ���   蔞����   ��ƃ�   ƃ�    ƃ�    �r������F�F ݕ�  ݕ�  ���  ݕ�  ǅ�      ݕ�  ݕ�  ݝ�  �/���_^ƅ8   ][��0�V�t$WV���b�����@  V�������t>h��h��h+  h���� ���N�O�V�W�F�G�N�O�V���W_��^� ����������̋T$SV��L$���ĉ�L$,�P�T$0�H�L$4�P�T$8�H�ΉP�W����؍D$P���������@  �P��D  �H��H  �P��L  �H��P  �P��T  ^��[� �������������j�hXd�    P��\�  3ĉD$XSUVW�  3�P�D$pd�    ��$�   j ��h;�  ����? �؄��h  ��P V���҅�������  ���H  ���B  ����g ��t\����g ��|Pj h;�  ���? �؄��  W���PQ j h���Ί��p? ��t���5�  ��u2ۋ��(�  ����  ����  j h;�  ���:? �؄���  V���  �4����Ί����  ����  ����  j h;�  ����> �؄��~  �D$DP�������L$DQ��蛟  �Ί���  ���S  ���M  ��l  Rh;	 ����> �؄��0  ���n�  ���  j h;�  ���> �؄��	  V��p  �r����Ί��9�  ����  ����  ���  Ph; ����E> �؄���  ����  ����  ���  Qh; ����> �؄���  �����  ����  ���  Rh; �����= �؄��l  ����  ���[  j h;�  ����= �؄��E  ��X  P���<�  �Ί��s�  ���$  ���  j h;�  ���= �؄��  V���  ������Ί��6�  ����  ����  j h;�  ���H= �؄���  ��   U�����  �Ί����  ����  ����  ���0e ��|1j hK�  ����< �؄��~  V��������Ί���  ���c  ���]  ����d ������)  j h;�  ���< �؄��2  jj���<�  �؄���   ���  Q���d�  �؄���   ݇�  �����$��  �؄���   ݇�  �����$�ʜ  �؄���   3��T$\R�ΉD$`�D$d�D$h�D$l��  �؄�t{�L$�CT �D$P���D$|    ��  �؄�tK��\  Q��軜  �؄�t7V���  ������؄�t%��8  R�����  �؄�t��(  W����  �؍L$�l$x�qT ���j�  ��t��tj U���; �؄�t���K�  ��u2ۊËL$pd�    Y_^][�L$X3���� ��h� ��j�h�d�    P��   �  3ĉ�$�   SUVW�  3�P��$�   d�    ��$�   3��l$$�l$�l$ ���������������D$0����L$4����T$8����D$ �D$ �D$<�L$@�T$D��I �D$P�L$(Q����  �؄��R  �D$$=;�  ��   ��   =;�  w~t`=;�  tF=;�  t=;�  ��  W���  ��������  ��B$W���Ѕ��Ä���  �D$��  W���  ��������  ��   Q���ٌ  ��Ɔ$  �  =K�  tG=;�  t =;�  ��  ��X  R��褌  ���n  �D$0P��聈  �؄��X  �D$�N  W��   �������;  W��p  �.������(  =; ���  ��  =;�  tE=;�  t/=; ���  �L$L$ t����  ��  2����  ��  V���3 ����  �T$R�D$0P�ωl$4�l$ �ѝ  �؄���  �   9D$,��  9D$��  ���a ���  ���w� =�o��m  �L$(Q�ωl$,蜆  �؄��S  �T$(R蘒 ���  �����  P����  �؄��(  ���  Q����  �؄��  ��$�   R���`�  �؄���   �L$H�}P �D$HP�ω�$�   �
�  �؄�u�L$HǄ$�   ������P �   �|$|���\  Q����  �؄�t�W���  ������؄�t��|$|���8  R����  �؄�t��|$|���(  P���^�  ��놋L$L$ t
����  �G2����  �==; �t =;	 �u/�D$P�D$,�� ����l  ��T$T$ t��2����  ����  ��u2ۃ|$$�t��������|$ tZ�|$ tS�L$0�,����tF��@  �����u7�L$0�T$4���ĉ�L$P�P�T$T�H�L$X�P�T$\�H�ΉP�$����A�D$xP���������@  �P��D  �H��H  �P��L  �H��P  �P��T  �Ë�$�   d�    Y_^][��$�   3��� �Ĝ   � �����j�h�d�    PQV�  3�P�D$d�    ��t$���   �D$   �%������   �D$�����N|�D$ �����Nx�D$����������L$d�    Y^������������V������V�V�N �T$�F    �T$�$�������T$��N8�\$�$�������T$�NP�\$���$����`/�Fh�d/�Nl�h/�Vp�l/�Nx�Ft�X����N|�P������   �E������   ^�9�����������̃�VW���D����|$3��D$�D$�D$P�L$Qh � @���`�  ��u_^��� �|$S�Ä���   V���[�  �؄���   �VR���F�  �؄���   �FP���1�  �؄���   �N Q���l�  �؄���   �V8R���W�  �؄���   �FPP���B�  �؄�to�|$|h�NQ���J�  �؄�tW�VhR���Y�  �؄�tF�FxP����  �؄�t5�N|Q����  �؄�t$���   R����  �؄�t�Ƅ   V���߆  �؋��f�  ��u2ۊ�[_^��� �����V�t$Wjj��h � @���84 ��u_^� �S�����$�?�  �؄���   �G�����$�%�  �؄���   �G�����$��  �؄���   �G P���6�  �؄���   �O8Q���!�  �؄�ty�WPR����  �؄�th�GP����  �؄�tW�OhQ�����  �؄�tF�WxR��譕  �؄�t5�G|P��蜕  �؄�t$���   Q��舕  �؄�t�Ǆ   W���t�  �؋�諼  ��u2ۊ�[_^� ������������̃�U�l$V3�W��D$�D$�D$P�L$Q�~h � @��� �   ���  ��u	_^]��� �|$S�Ä�t3V��覎  �؄�t%W���8�  �؄�t�? u���fZ ��|�   ��蔾  ��u2ۊ�[_^]��� ��VW�|$j j��h � @���h2 ��u_^� �SP����  �؄�t"�v��u����Y ��|�   V��譐  �؋�蔻  ��u2ۊ�[_^� ������QU�l$�������D$P���D$    �o  ��tF�L$��~>SV��Qj覭���L$����VQ���$�  �؄�tV��������t	V蜭����^��[]Y��̃�X�L$@�d���L$(�[���L$�R���D$@P����  ����   �L$(Q����  ��t�T$R���  ��to�D$P���R  ��t_�$Q���~  ��tPS�T$R���~  �؄�t:�D$P�L$0Q�T$LR����� �D$�D$ݗ�   �L$ݟ�   ���   ���   ��[��X������������U������|S�L$P����D$ P���1~  �؄��v  �L$$Q���~  �؄��`  �T$PR����~  �؄��J  �D$HP���~  �؄��4  �L$@Q���i~  �؄��  �T$8R���S~  �؄��  �D$0P���=~  �؄���   �L$(Q���'~  �؄���   ���D$(���������A{	������Az����'�T$(���D$0��������A{������Az������Xe�T$0��Wjdjd��(�\$ 3��|$T�\$��$�   �D$l���\$�D$t�\$�D$|�$R��P�U�����<�L$hQ���F������@  �H��D  �P��H  �H��L  �P��P  �@��T  ��[��]����������̃�SU�l$VW�͋��|����D$P�L$Q����  �؄���   �D$=  �wgtG-  t+��t����   ���  �$������   ����������u��X  R�����������`�D$D$t
����  �L2����  �B=  �t%=	  �u4�L$L$t
����  � 2����  ��T$T$t��2����  ���6�  ��u2ۃ|$�t������_^]��[���������̃�SU�l$VW���   芊����    �hY���ݕ�   ݝ�   ǅ�   F   ǅ�      ƅ�   �I �t$�D$P�L$$Q���k�  �؄�tD�D$ -  t��u�����������   P���n������؋��r�  ��u2ۃ|$ �t��u�_^]��[���������̃�dSU�l$pVW�͋��������T$�\$$���D$P�L$Q�����  �؄���  �D$=  �|  �i  �������Z  �$�`��T$R����z  ���@  �D$$P����z  ���-  ��X  Q�����������  ���  �������  �����������  ��p  R���z  ���  P���z  ��x  Q���sz  ���  R���ez  ���  �L$\�����L$D�����L$,�����D$\P���z  �؄�t �L$DQ���uz  �؄�t�T$,R���cz  �؍D$,P�L$HQ�T$dR���  �� ���G  ��  P����y  �؄��/  ��  Q����y  �؄��  ��  R������������   �D$  ���   =	  ���   tv=  tZ=  �t/=  ���   �D$D$t����  �   2����  �   �L$L$t����  �   2����  �   ��   R������������o�D$D$t
����  �[2����  �Q=  �t6=  �uC�D$�L$���t��u0��u,ǅl     � ǅl     ��D$D$t
ǅ�     ��葶  ��u2ۃ|$�t���L���_^]��[��dË��5�#�8�8�8�8�8�8�C�������������������j��览  ���
wM�$�H��   �A�   �:�   �3�   �,�   �%�   ��   ��   ��	   �	�
   �3Ʉ�tDQ���E�  ��t8�G�����$�щ  ��t$�G(�����$轉  ��t�G �����$詉  ����������������������������������̋D$�T$��    +����QR�B������ ������������VW�|$��;~tzS3�;�~Y9~~�~�N��PWQ����;ÉFtO�V;�~,U��+ʍ,�    +����    �U+ʍ�SR�� ��][�~_^� �F;�t�SP�B�Љ^�^�^[_^� ����SW�|$����~uU�l$��|kV�t$��|a;�t]�C�/;�S;�O�K�>;�~�;�}��P���&����C��    +����R��    +͍ȍ�    R+΍�R�d� ��^]_[� ���������̋Q2���t(�I��~!V�t$��t��~Vh�   QR��: ���^� �����������̋Q2���t(�I��~!V�t$��t��~Vh�   QR�: ���^� �����������̋D$�L$����PQ�{������ ����̋Q2���t(�I��~!V�t$��t��~Vh(  QR�E: ���^� �����������̋Q2���t(�I��~!V�t$��t��~Vh(  QR��9 ���^� �����������̋D$�L$i�(  PQ�ۢ����� ����̋Q2���t%�I��~V�t$��t��~VjLQR�9 ���^� ��������������̋Q2���t%�I��~V�t$��t��~VjLQR�X9 ���^� ��������������̋D$�L$k�LPQ�>������ �������̋D$S��VW��    ���݀�   ݛ�   ݀�   ݛ�   ���   ���   ���   ���   ���   �   ���   P���   ����_^��[� �������SU�l$��VW�    �����݅�   ݛ�   ݅�   ݛ�   ���   P���   衉�����   ���   ���   _���   ���   ^���   ]��[� ����j�h�d�    PQ�  3�P�D$d�    �L$�L$���D$    t�6@ �L$d�    Y��� ����j�h��d�    PQV�  3�P�D$d�    ��t$�NH�D$	   �H����ND�D$�;����N@�D$�.����N<�D$�!����N8�D$�����N4�D$�����N0�D$������N,�D$�����N(�D$������N$�D$ �Ӏ���N �D$�����À���L$d�    Y^�����VW�|$��;�t4��O��GQ�^�N�.����G�^�G �^ �G(�^(�W0�V0�G4�F4_��^� ��������̃�V���@WWtJ�@W��HWhPW�^�N�ԇ���XW�^�`W�^ �hW�^(�pW�N0�tW�V4�|$�D$P���D$    ��p  ����   �L$�����c��   �T$R���D$    �p  ��t8�D$P��r ���NQ�ω�%q  ��t�V R���q  ��t�F(P���q  �|$e|o���D$    t+�L$Q���Xp  ��t�T$R�y �F0���F4P���9p  �N4��|��~�F4   �|$f|��t�NQ���p  ��t��V����t  _^��� ���������j�hˀd�    PQV�  3�P�D$d�    ��t$�Nd������D$    �����ƋL$d�    Y^�����������������j�h�d�    PQUVW�  3�P�D$d�    ��l$�� ���   ���D$    �<�����D$�P~����    �hY���ݕ�   ݝ�   ǅ�   F   ǅ�      ƅ�   �ŋL$d�    Y_^]�������j�hF�d�    PQSUVW�  3�P�D$d�    ��l$� � ���   ���D$     �~����    �hY���ݕ�   ݝ�   ���D$ �}��ƅ�   ƅ�    ƅ�    �ŋL$d�    Y_^][�����������j�hx�d�    PQV�  3�P�D$d�    ��t$�~�����D$    �$}���F�F �ƋL$d�    Y^������������j�h��d�    PQVW�  3�P�D$d�    ��t$�~8���}�����V���V�D$    �V�    �V �V(�^0�|���ƋL$d�    Y_^���U�������   SV��W��X  ��~�����D$4u�D$4�7���͛���L$h��������$�   ������$�   �z�����$�   �n�����$�   �b���P��$�   �U���P��$�   �H���P�L$t�>���P�������؍D$XP��$�   Q��$�   R��$�   P��$�   Q�T$tR��貝�����L$PQ�D$L�T$<R�D$DP�L$PQ�T$\R�D$hP��������ȋǃ��L$@t��t�,1��`���T��T$4�}PRh,�W� �����~ ����   ݄$�   ��`�\$X݄$  �\$P݄$   �\$H݄$@  �\$@݄$8  �\$8݄$0  �\$0݄$(  �\$(݄$   �\$ ݄$  �\$݄$�   �\$݄$�   �\$݄$�   �$h��W�i~ ��h��$�   P�������L$hQ��$�   �f��݄$�   �� �\$݄$  �\$݄$  �\$�$h��W�~ ��(�|$H tO�D$X��0�\$(݄$�   �\$ ݄$�   �\$݄$�   �\$݄$�   �\$݄$�   �$h8�W�} ��8�|$@ t,�T$P�D$8�L$<R�T$HP�D$TQ�L$`RPQh��W�} �� ݆�  �� ��'�����\$݆�  ���\$݆x  ���\$܎p  �$h8�W�E} ��(����| _^[��]� ��j�h�d�    PQV�  3�P�D$d�    ��t$�N �����N8�����NP�����Nx�z���N|�D$    �z�����   �D$��y�����   �D$��y�����D$�����ƋL$d�    Y^�����������̃�V����@W�D$    �D$    tJ�@W��HWhPW�^�N�E����XW�^�`W�^ �hW�^(�pW�N0�tW�V4�D$P���\i  ��t�L$Q���Li  �L$��
wW�$����   �N�   �F�   �>�   �6�   �.�   �&�   ��   ��	   ��
   ��    ��t)�VR���gi  ��t�F(P���Xi  ��t�� V���Ii  ^���d���$�,�4�<�D�L�T�\���������QSUV�t$W�����B ����   ���   ��   j h5�  ���j �؄���  j j����~  �؄�t���  P���!y  �؄��D$    t+3퐋D$;��  }���  �V�2 �D$�؃�L��u؋��ѣ  ���q  ���k  j h1�  ���� �؄��S  V���   �}����Ί�蔣  ���4  ���.  j h2�  ��� �؄��  V��  �P����Ί��W�  ����  ����  j h3�  ���i �؄���  V���  �����Ί���  ����  ����  j h4�  ���, �؄���  V��P  �����Ί��ݢ  ���}  ���w  j h5�  ���� �؄��_  ���  U�Ήl$�w  ����D$    ~Q3�I ��tHj h;�  ��� �؄�t���  �V�����Ί��a�  ��u2ۋD$���Š   ;D$�D$|����=�  ����  ����  j h6�  ���O �؄���  ���  U���w  ����D$    ~W�D$    ���tJj h;�  ��� �؄�t���  L$V������Ί�迡  ��u2ۋD$�D$(  ��;ŉD$|���蛡  ���;  ���5  j h7�  ��� �؄��  ���  U�Ήl$�qv  ����D$    ~O3퐄�tHj h;�  ���n �؄�t���  �V�*����Ί��!�  ��u2ۋD$����(  ;D$�D$|������  ����  ����  ���  Qh8  ����
 �Ί��Ѡ  ���q  ���k  j h9�  ���� �؄��S  ���  R���u  �؄ۋ�   t
P���u  �؋��~�  ���  ���  j h:�  ��� �؄��   ��  P���w  �؄ۋ�  t
P���Du  �؋��+�  ����  ����  ��$  Qh<  ����8 �؄���  �����  ����  j h=�  ��� �؄���  V��(  �K����Ί��  ���b  ���\  j h?�  ���� �؄��D  V���  �~����Ί�腟  ���%  ���  ���~s����~1j h1�  ��� �؄���  W���
x  �Ί��A�  ����  ����  ��  Rh2 ����N �Ί���  ����  ����  ��   Ph3 ����" �Ί���  ����  ����  ���"= ���Q  j h4�  ���� �؄��[  jj���vy  ݇�  �����$�Cu  �؄��  ��  Q���;u  �؄���   ��  R���ss  �؄���   ��  P���[s  �؄���   ��  Q���Cs  �؄���   j jh � @��� �؄���   V���   �����Ί����  ��u2��o��tk���  R����t  �؄�tW�GP���t  �؄�tFV�O � ����؄�t7���  ���  Q�����  �؄�tV�������؄�tV���  �u����؋��|�  ��t ��tj j���� �؄�t���\�  ��u2�_^]��[Y� ������������V�t$W�����; ��u7Sj h  ���M �؄�t�Ǩ   �l����Ί���  ��u2ۊ�[_^� V���}���_^� ��������V��~ ���t%�F��tj P����F    �F    �F    ^�����������VW�|$��;�tJ�G��_�F    ��^� 9F}P������N��t#�G��    +���҉F�GRPQ轸 ��_��^� ���V��L$��|<�F;�}5+���P�APQ�������F��F�V��    j8+ȍ�j P�\� ��^� �����V��~ ���t%�F��tj P����F    �F    �F    �D$t	V��u������^� ������SVW�|$W��������(  �@��(  ��(  R�Њ�8  ��8  ��@  ��@  ��D  ��D  ��H  ��H  ��L  ��L  ��P  ��P  ��T  ��X  ��T  R��X  ��u����\  ��\  ��`  ��`  ��d  ��d  ��h  ��h  ��l  ��l  ��p  ��p  ;�t"� ��@�Y�@�Y�@�Y�P �Q �@$�A$���  ���  ���  ���  ݇�  ݞ�  ���  ݇�  Pݞ�  ���  ݇�  ݞ�  ݇�  ݞ�  ݇�  ݞ�  ݇�  ݞ�  ��t�����  Q���  �������  ���  ���  ���  ���  ���  ���  R���  �������   ��   W���t���G�C�O_��^�K[� ���������������j�h1�d�    PQ�  3�P�D$d�    �L$�L$���D$    t������L$d�    Y��� ����j�h��d�    PQSV�  3�P�D$d�    ��t$����3ۉ\$ǆ(  ����,  ��0  ��4  ��@  �D$�`�����X  ��l����ݖp  ���  ���D$ݖx  ���  ݞ�  ���  ���  ���  ���  ݞ�  ��������  �D$�������  �D$������   �D$�;������D$�o����ƋL$d�    Y^[��������������j�h�d�    PQSVW�  3�P�D$d�    ���|$��   �D$   �3k�����  �D$�S������  �D$�������  �D$�k����X  �D$��j��3�9�4  ��(  �\$���t�F;�tSP������^�^�^���D$������~���L$d�    Y_^[����������������j�hY�d�    P��SUVW�  3�P�D$d�    �ًk���|   �|� ���d$ �s��t$���   �D$$    �4j�����D$$�����& �Ch�   �j P�S� �K��ωL$�L$�D$$   t�T�������   ���D$$����}��C    �L$d�    Y_^][�������SUVW�|$����}V3�9n�  �~��x%�������    �N����������   ;�}�N��PUQ����_�n�n�n^][� �F;�}n�N��PWQ����3�;ŉF��   �V��+ʍ�����Q���UR�\� �F��;�}"������+�F�P���+����à   ��u�~_^][� ~Q���;�|"��+�������N��6�����   ��u�9~~�~��F�RWP�Ή~��3�;ŉFu�n�n_^][� ������������UW��3�9o� �t:V�w��xS�����O��Ž������   ;�}�[�O��PUQ���҉o^�o�o_]�������������V�������D$t	V�o������^� ��V��F�V����;�uJ��   v��|��� ;�}�������   ��;�}8P��������N����F���N^�N�����F����V��R�����N����F���N^����j�h��d�    P��   SUVW�  3�P��$�   d�    ��F�n;ŋ�$�   ��   ������   v��|��� ;�}�ȍ<����   ~�< �F��tx��+ȸgfff���������xa;�}]�L$�1���S�L$Ǆ$�       ����9~}W��������F����N�T$��R�F������L$Ǆ$�   ���������$;�}W�������F����N��S�F������$�   d�    Y_^][�Ĭ   � �������������SUVW�|$����}S3�9n��   �~��x"��k�L���$    �N��v�������L;�}�N��PUQ����_�n�n�n^][� �F;�}f�N��PWQ����3�;ŉF��   �N��+�k�Lk�LR�UQ�ժ �F��;�} �؋�k�L+���F�P��������L��u�~_^][� ~M���;�|��+�k�L����N��������L��u�9~~�~��F�RWP�Ή~��3�;ŉFu�n�n_^][� �����������UV��3�9n�(�t6W�~��xS��k�L�N��V�������L;�}�[�N��PUQ���҉n_�n�n^]�V�������D$t	V�k������^� ��j�h��d�    P��SVW�  3�P�D$d�    ���_��x`��i�(  ���    �O�������Gh(  �j P�t� �O��ΉL$�L$�D$     t��������(  ���D$ ����}��G    �L$d�    Y_^[���������V��N�V;�uL��k�L=   v��|��� ;�}�������   ~�	;�}7P���j����N��k�LF���N^�k�LN������Nk�LNQ�������N��k�LF���N^���������UW��3�9ot<V�w��x!S��k�L��    �O���������L;�}�[�O��PUQ���҉o^�o�o_]�U������4SVW����b������T$�T$�N�$������N ��������   ��@WtJ�@W��HWhPW�_�O�Bj���XW�_�`W�_ �hW�_(�pW�O0�tW�W4���   ��@WtJ�@W��HWhPW�_�O��i���XW�_�`W�_ �hW�_(�pW�O0�tW�W4��  袛�����  藛��3ۿ   ���  ���  ���  �i�����P  農�����  �C������  �8������  �-����`/���  �d/���  �h/S���  �l/SS��  ���  ���  ��  ��   ǆ�  ������   �M��j��L$@��  ǆ  ������  ��J���L$<��  ��(  ��  ��$  �ͫ����ݖ�  ǆ�  F   ݖ�  ǆ�     ���  ���  ���  ݞ�  ���  ����_^[��]��UV��3�9n��t<W�~��x!S��i�(  �N��3�������(  ;�}�[�N��PUQ���҉n_�n�n^]�����������V�������D$t	V�[g������^� ��j�h��d�    PQSV�  3�P�D$d�    ��t$�a��3ۍN�\$�T����N �������   �D$�l������   �D$�\�����  �D$�������  �D$�|������  �D$�l�����P  �D$����ǆ�   ����  ���  ���  �����  ���  ���  ���  ���  ���  ���  ���  ��  �D$
��H����  ��H����(  �Ū����ݖ�  �   ݞ�  ǆ�  F   ǆ�     ���  ���  ���  ǆ�  (����  ���  ���  ���D$���  ���  ������ƋL$d�    Y^[�������j�hO�d�    PQV�  3�P�D$d�    ��t$���  �D$   �u�����(  �D$
�e������  �D$	�������  �D$�u������  �D$�������  �D$�%^�����  �D$�� ���  �D$�� ��  �D$�� ���   �D$��]�����   �D$��]���N �D$ �h������D$�����]���L$d�    Y^�����������j�h{�d�    P��,  �  3ĉ�$(  SUVW�  3�P��$@  d�    ��$P  ��F�n;���   ��i�(  ��   v��|��� ;�}�ȍ<����   ~�< �F��t|��+ȸ�=`������
�����xc;�}_�L$�o���S�L$Ǆ$L      ����9~}W������F��i�(  N�T$��R�F������L$Ǆ$H  �����+����&;�}W���]���F��i�(  N��S�F������$@  d�    Y_^][��$(  3��� ��8  � ���������j�hхd�    P��	  �  3ĉ�$ 	  SVW�  3�P��$	  d�    ��$$	  ��P���2��҉D$��Pj ���҄��\  �D$P�L$Q�����  ���C  �D$�������"  ��0��$����$�   �������$�   P��Ǆ$ 	      ��������t��$�   Q���  �������$�   Ǆ$	  ����������   �L$ ������T$ RWǄ$$	     ��������t�D$ P���  �����L$ Ǆ$	  �����h����h��$�  ��h�����$�  Q��Ǆ$ 	     ��������t��$�  R���  ������$�  Ǆ$	  �����-�������   ����������  ��������L$��PQ���ҊË�$	  d�    Y_^[��$ 	  3��� ��	  � ���j������� ��̃�p�  3ĉD$lSUV��$�   ��W�l$,��l$,�D$P�L$43�Q�Ή|$8�|$�|$ ��  �؄���  �D$0=1�  �  �
  ��߃���  �$�l����   V���:���W���   ��������]  V��  �K������J  V���  �8������7  V��P  蕪�����$  �Ÿ  �������T$@R�Ή|$<�|$P�|$T�J  9|$@����  ����  �D$LP�L$<Q���4�  �؄�t,�|$8;�  t2���������V��衯���؋��H�  ��u2ۃ�;|$@|��  ���  ���'����T$4R�Ή|$H�|$`�|$d�I  9|$4���i  �I ���^  �D$\P�L$HQ��觑  �؄�t,�|$D;�  t2�������V�������؋�軇  ��u2ۃ�;|$4|��  �l$,���  �������T$(R�Ή|$@�|$X�|$\��H  �؋D$(P�����9|$(��  ��    ����  �L$TQ�T$@R����  �؄�t,�|$<;�  t2��������V���t����؋���  ��u2ۃ�;|$(|��m  �|$�b  9|$�X  �D$dPj����>  ���C  ���  Q�Ή|$�KH  �؄��'  �T$R���5H  �؄��  �D$P�AS ����   ��  ��  Q�Ή|$�H  �؄���  �T$R����G  �؄���  �D$P�R ����  �  V��(  �=������  V���  �������  U���L  ���z  =<  ���  ��  =4�  ��   =5�  tG=8  ��L  �T$�D$�ʃ��;�wr��   �w���  �$  h��h��h`  �  �L$Q�T$$R�Ή|$(�|$$�|$��]  �؄���  �|$ ��  9|$��  �D$P����F  9|$����  ����  ;|$��  �L$,V���  ��������� �؃���u��  �L$Q�T$ R�Ή|$$�|$�f]  �؄��b  �   9|$�S  ���  P����F  �؄��;  ��  Q����F  �؄��#  �T$$R���1F  �؄��  �D$$P��P ����  Q�Ή�  �F  �؄���  �T$$R����E  �؄���  �D$$P��P ��9|$��  ��  �L$ Q�T$LRh � @�Ή|$T�|$,��  �؄�tV���   �I����Ί���  ��u2ۃ|$�e  ���  P���G  �؄��M  �|$�B  �MQ���1F  �؄��-  V�M �����؄��  �|$�  ���  W���{S  �؄���   �|$��   V���^����؄���   �|$��   V���  轓���   �T$�D$�ʃ��;�wr��  �w��$  �   h8�h��h�  �x=2 �t==3 �uw�T$�D$�ʃ��;�wr��   �w��   �Rh��h��hw  �4�T$�D$�ʃ��;�wr��   �w��  �hp�h��hk  h���ͳ ����蓂  ��u2ۃ|$0�t�������L$|_^]��[3�藓 ��p� �I �����������)�6���=�6�6���������������VW�������|$���� ��W��u
�O���_^� �e���_^� �A+A���������̋D$�L$VW�   ��;u��������s��t^��8+�uE��������tG��8+�u.��������t0��8+�u��������t�� +�t�Ҹ   _���^�3�_^�����̃�V��F;F��   U3�;���   3�9nW�n�D$�l$~i�l$S�D$�~�8Shp/�$������u,�L$;L$~��/�C�D/�K�L/�S�T/�D$���D$�D$��;F�D$|��D$3�[;F}D;ŉF~:�   ;ǉ~~1�F�N���P���P�m������~�V;V|�_]^��Én_]^����������3��A�A�A������k��������������V�t$W�|$VW�O�������u��V��W�;�����_^�����̋D$�L$�@���PQ�p����� �̋T$�A�IR�T$R�T$RPjQj j� �� � �������̋T$�A�IRPjQj j�X� ��� �̋T$�A�IR�T$RPjQ�7� ��� �V��F9F|�~ ~l�N��t#��~�����t��~h��jPQ�H ���~ ~/S�^W�~�����L�Qhp/��"������t
������~�_[�V�F    �V^��V��FW3�;F~�m����F��~9Fu9~u�F_^Ë�_^��VW�|$j j��h � @����  ��t4�|$ ��t�&�����O���SV���y  �ϊ���{  ��u[_^� ��[_^� ����������̃�SV3���W�|$�F�F�F�D$�D$�D$P�L$Qh � @���+�  �؄�t"�|$t2��
V����K  �؋��~  ��u2ۀ|$ ��t����_^��[��� ����_^��[��� ����������QW���G+G��� ~�F����G��~g�O�T$h��jPQR�ۭ �����D$u^S�_V�w;�}PU�o�������$    �D$WP��������t$����;�|�D$]^[_Y� �D$    �D$������]^[_Y� ����������̋D$9A}	�D$�*��� ����������̃�$�  3ĉD$ V��F;F��   �N��t#��~�����t��~h��j PQ�� ���~ ��   �t/�x/3��~ �D$�D$�D$�D$�D$�D$�D$�D$ �p/W�=|/�D$�L$�T$�|$�D$�L$�T$ �|$$~DU�nS�^�����|(��L$WQ�c�������u���T$ WR�N�������u
����ۉ^�[]�F    _�F�F�L$$^3��+� ��$�������������̃��  3ĉD$V��F;F��   �N��t#��~�����t��~h��jPQ� ���~ vr�L$�z   �~ �p/�t/�x/�D$�|/�L$�T$�D$�D$    ~.S�^W��~���T��R�D$P�k�������u
������~�_[�F    �N�N�L$^3��I� ��������������QW���G+G��w� v�����G��v_�O�T$h��jPQR�� �����D$uUU�oV�w;�}G���S���L$SQ���������t$����;�|�D$[^]_Y� �D$    �D$봍���[^]_Y� ����V��~ ��t%�F��tj P�$��F    �F    �F    ^�����������VW�|$��;�tD�G��_�F    ��^� 9F}P脚���N��t�G�F�W�@���PRQ�Ó ��_��^� ��������̋D$V��3�;���$�N�N�N~P���ܝ����^� ������V��~ ��t%�F��tj P�$��F    �F    �F    �D$t	V��P������^� ������V��~ �,�t%�F��tj P�8��F    �F    �F    �D$t	V�P������^� �����̋�3ɉH�H�H� @�������������̋D$V��3�;��lI�N�N�N~P����s�����@�^� 3�V��F�F�F�D$P�lI�pI�@���^� ����̋D$V��;�tP�Ϡ����^� ��������̋�3ɉH�H�H� T�������������̋D$V��3�;���$�N�N�N~P���L������T�^� 3�V��F�F�F�D$P��$��$�T���^� ����̋T$�A�IVR�T$�rVRPjQj j� �� ^� ������̋D$V��;�tP�_�����^� ��������̋�3ɉH�H�H� h�������������̋D$V��3�;���I�N�N�N~P���ܕ�����h�^� �D$V��;�tP�_�����^� ��������̋�3ɉH�H�H� |�������������̋D$V��3�;���H�N�N�N~P���������|�^� ��3ɉH�H�H� ��������������̋D$V��3�;���J�N�N�N~P��輕�������^� �D$V��;�tP��Q����^� ���������VW��3�j W��[�~�~�~��[;ǉFt:�N�� }�    +���R���WQ�� ���~�~_�F    �����^É~�~�~�~_�����^����������̋D$V��W3�;���[�~�~�~~P��p���~�~_�����^� ����������V��W3�9~�~�~��[t�F;�tWP��[�~�~�~_^���������������VW�|$��;�tW讝���G�F�O�N_��^� �����������VW�|$j j��h � @����  ��t&S������V���to  �ϊ��kr  ��u[_^� ��[_^� ��������̋D$jP�d���� ̃��  3ĉD$�D$�T$�$�D$ �D$�T$�T$$�$P�T$�����L$���3���賅 ��� ���VW��3�j W����~�~�~���;ǉFt?�V�� }�    +ʍ���Q����WP�� ���~�~_�F    �����^É~�~�~�~_�����^������V��W3�9~�~�~���t�F;�tWP����~�~�~_^��������������̃��  3ĉD$�D$�T$�$�D$ V�t$,�D$�T$�T$(�D$P�T$�t�����t	��t�H��L$3҅���^3̊�茄 ��� ������������VW��3�j W�,��~�~�~�8�;ǉFt:�N�� }�    +���R���WQ�܈ ���~�~_�F    �����^É~�~�~�~_�����^�����������V��W3�9~�~�~�,�t�F;�tWP�8��~�~�~_^���������������VW�|$��;�tW�~  �G�F�O�N_��^� �����������V��~ �lIt%�F��tj P�xI�F    �F    �F    �D$t	V�I������^� ������V��~ ��$t%�F��tj P��$�F    �F    �F    �D$t	V�_I������^� ������j�h�d�    PQVW�  3�P�D$d�    ���D$    �t$ ���D$    �P� �G�j �NQVPjWj j�D$8    �D$,   � �� �ƋL$d�    Y_^��� �������������V��~ ��Ht%�F��tj P��H�F    �F    �F    �D$t	V�H������^� ������V��W3�9~�~�~��[t�F;�tWP��[�~�~�~�D$t	V�4H����_��^� ���������̃��  3ĉD$�|$( �T$S�\$(VW�|$,��L$$�L$�T$�|$�\$tB���ĉ�P�x�ΉX�o������Ä�t�D$P����{���L$_^��[3��D� ��� ���V��W3�9~�~�~���t�F;�tWP����~�~�~�D$t	V�dG����_��^� ���������̃��  3ĉD$�|$0 S�\$(U�l$(VW�|$,��L$8�|$�l$�\$�L$ tSj ���ĉ8�h�X�H�������������D$tU�D$Php/� ������t2�_^][�L$3��b� ��� �D$�̋��T���L$ �T$<�8�h�X�H�P�D$�L$$_^][3��%� ��� �����V��W3�9~�~�~�,�t�F;�tWP�8��~�~�~�D$t	V�DF����_��^� ����������QSUV��F+FW�|$�_�9G�\$}P���i��3�9n~73ۋF�<Whp/�������u
�L$W�z������;n|Ӌ\$�|$�G_^]+�[Y� ��������������Q�L$���$    t,�9 t'�D$��t�8 tPQ�D$P�#� �����$t��u3�YËD$��t	�D$�® ��������������̋T$�D$�ʁ�   ��� ��wr���w���h �h��hM  h��贞 ���    2���������̃|$ w�D$r���w���h<�h,�h[  h���p� ���    2�����̃�(�  3ĉD$$U�l$0��V�t$@W�|$@t%~��t��u_�D$ �D$^]�L$$3��~ ��(�S�\$@�Ã��D$�<  ����   ��tZ�C���wH���C  ��$    ����~)S�L$WQ�}� ����ۋ�t���T�������u���u��  �D$ ��   ����   ��I ��O���W���_���\$�_���\$�_���\$�_���\$�_��\$�^�\$�����^�\$���^�\$�����������������������s����]��tY��O���W���_��������������������u��%��t!��I ��O��������������u�L$4�D$[_^]3��| ��(��������������SV�t$��W�|$��w�����v0��$    ��Ph������҄�t/��  ������w�r�����wׅ�w��v��PW����_^[� _^2�[� _^�[� ���������������SV�t$��W�|$��w�����v0��$    ��Ph  ����҄�t1��  ������w�r�����wׅ�w��v��P��W����_^[� _^2�[� _^�[� ������������̊�x@  $�������̋�x@  ��$������j�hH�d�    P�  3�P�D$d�    �D$P���   �D$    �(B���L$�D$�����w:���L$d�    Y��� ����̅�u2��V�ph�/V�j������u^h�/V�X������uLh��V�F������u:h�/V�4������u(h 0V�"������uh��V�������u2�^ð^�̋A���Шt�A�I��|	��r���3�3�������������̃|$ ��@  ��@  � ��������̊�@  ���������̃|$ ���@  ���@  � ��������̊��@  ���������̃|$ ��|@  ��|@  � ��������̸2   ����������̋L$������3�����   �$��	�   � �   � �   � �   � �   � �   � �   � �   � �	   � �
   � �   � �   � �   � �   � �   � �   � |	�	�	�	\	d	l	�	�	�	�	�	�	�	�	�	�	�	�	�	�	t	�	��������;�s2+ȃ�|+��t#�|$ t�H�
��J�����
�H�J���3���������;�sN+Ѓ�|G��t?�|$ t�P��P�Q�P�Q��Q������P�Q�P�Q�P�Q���3�������������;���   +Ѓ�|��tw�|$ t:�P��P�Q�P�Q�P�Q�P�Q�P�Q�P�Q��Q������P�Q�P�Q�P�Q�P�Q�P�Q�P�Q�P�Q���3�����������������Q3҅���;��$sN+ȃ�|G�|$ t�H�P�$�H�T$����P�$�H�T$�P���T$�L$t94$t3�Y���������������̃|$u�L$�������Q�L$�t�������t��t�L$��F    �����������̃�V��;�W�|$�D$    �D$    �D$    sw+ȃ�|pW�L$����������t_W�T$�����������tLW�T$����������t9;�s3+���|,�T$f�L$�f�T$f�Kf�S��K�P_�S��^���3�_^������������̃�(�  3ĉD$$�D$4S�\$0V�t$@�L$S���x�������u^[�L$$3���u ��(Ã���|$8U�L$�L$S��u�L$�����t$ ����L$�/���������  3����l$�}  ���u  ���k  �|$D��  u�T$<3Ƀ�1;�rw;�r�D$����D$ �9  ���1  S�\$$���n����؃����  �D$��tP�T$$R���������   �|$ t~�D$8P���  �ϋ��y���������   ����L$�L$�L$<Q�L$<�t$�������؃�����   �L$�ɋt$��   ����   ;���   ��+Ù;�|};�rwދT$8R�L$�׋������������tZ�D$ Pjj �e� �L$0QjP�X� �T$>RjP�K� �L$LQjP�>� ��03�9D$]��#�^��[�L$$3��t ��(ËL$0]^[3�3��t ��(������U�����x@  u�y uy�yus���@  ��tiS�\$��t_�; tZVW��3����  }J�> |E�N��|=��   5�F��t.�8 t)�< u#SP�3$ ����t�v����u�_^[��]� �._^[��]� ��������������j�h{�d�    PQV�  3�P�D$d�    ��t$�N�p���N�D$    ������ƋL$d�    Y^���������������̃�������������U���������S�KW����������z��F��������Au�V�F��������Au�V�F�^����������Au��F ��������Au���V ���F(��������Au���V(���F0�~0��������Au������F8��������Au�^8����F@����������Au�^@��؋��!���������W�D$SP�>�����VH�P�NH�Q�P�Q�P�Q�P�Q�@���A�������x _[��]���̸�W�����������j�h��d�    P��V�  3�P�D$d�    ��t$��� ���   �D$$    �t�舓���D$P��W�D$(�F(    � ����N�P�V�H�N�P�V�`/�F�d/�N�h/�V �l/�F$Ɔ�    �ƋL$d�    Y^�� �����������j�h�d�    PQV�  3�P�D$d�    ��t$�t����   �D$    ��� ���D$�����P� �L$d�    Y^�����������������̋L$h���8���   � ���������̋�t@  ���������̋A4������������̋D$��V��u3�^� ��RW�~�σ�P�D$�NP���҉~_3�^� ����������SV�t$3ۃ�|��~!��2|&�gfff������������+�u
�q^�[� h��h��h�3  h���Y跏 ��^��[� ������������̋��@  ��t�L$P�D$PjQ蕕 ��� 3�� ���������V�񋖘@  3���W��   ���@  ��tw���@  �|$�8;��@  r0��P���҄�u_3�^� ���@  �L$PWjQ�٣ ��_^� �T$WR�P�w ��@  ���@  ��;��@  v���@  ��_^� �D$�L$RPjQ荣 ��_^� �W�����@  �ɰtm���@  ��tc���@   vZSV���@  QVjR�P� ��;��Ä�t$���@  ;�t+�jP���@  P�� ����u2�^��Ǉ�@      Ǉ�@      [_���VW�����@  3���tPP�E� ����$|��sh��h`�h4  h���� ��������@   t0���@   v'��@  _��^�h4�h`�h$4  h���Ǎ ��_��^����������������QV�񋎘@  �ɰt\S2ۄ�x@  tNQ账 ����u(���@  Pj�L$jQ脓 ���@  R茦 ����t[�^YË��@  jj�P�� ����[^Y��SV��2ۃ��@   to���@   W�|$t ���@  �x;��@  w���@  _^�[� ��B�Ћ��@  jWQ荥 ����t�h��h��hi4  h���͌ ��_^��[� ^��[� �����������SV��2ۃ��@   tD��P�ҋD$���@  j PQ�'� ����u^�[� h0�h�h�4  h���`� ��^��[� �����̋�3ɉ�H�H�H�H��������������V��F��t�N�H�F��t�V�P�F��tP��J�����F    ^����������̋��@  ����������2����@   t/�T$��|��@  �� V���@  W����;�w
򉱤@  �_^� ���2����@   t�D$3�;��#Љ��@  �� �������������̋��@  ;��@  ���VW�|$����vH�T$��t@���@  ���@  ;�v+��3�;�v����v���@  W�PR��s ����@  ��_^� _3�^� �����3�� ����������̋T$��V��t0�N��t)�F��~"W�|$WjPQR�ɉ ����_t
+F^��� ���^� �������������̋A��~�I���D��3�������������VW�|$��;~tkS3�;�~J9~~�~�N��PWQ����;ÉFt@�N;�~��+�iɐ  iҐ  R�SQ��n ��[�~_^� �F;�t�SP�B�Љ^�^�^[_^� ���VW�|$��;~teS3�;�~D9~~�~�N��PWQ����;ÉFt:�N;�~��+���R���SQ�Tn ��[�~_^� �F;�t�SP�B�Љ^�^�^[_^� ���������j�h!�d�    PQ�  3�P�D$d�    �L$�L$���D$    t��Z �L$d�    Y��� ����j�hQ�d�    PQ�  3�P�D$d�    �L$�L$���D$    t�6)���L$d�    Y��� ����S�\$��VW�|$��w�����v9��Ph����҄�t!��  ����SW���%�����t_^�   [� _^3�[� ��PW��_^��[� �������������V��~ �l�t%�F��tj P�x��F    �F    �F    ^�����������VW�|$��;�t>�G��_�F    ��^� 9F}P�Tw���N��t�G�F��P�GPQ�p ��_��^� ���������������W����u2�_ËD$�@��Vt��2uG�wVh 0�%�������u-V��OQh�/��������t��Wh|����������t^�_�^2�_�������̅�u2��V��� ����tW���u�������u���w� ����u�2�^ð^���������̋A(��~�I$V��W�|$���t
�   �_^� �T$3ɉ
�J�J�J�J�J�J�J� �����������V��~ �l�t%�F��tj P�x��F    �F    �F    �D$t	V��,������^� �����́�  �  3ĉ�$�  ��$�  ��$�  SV��$�  ��$�   ��$�  ��$�   ���$�   ��$�   �B3�W�Ήt$0�\$�Ћ�$�  ��$�  3�;ӉD$|w;�v
;�rwa;�s]��t@  ��$�  ��$�  �D$3Ƀ~2�\$D��=  ��   �L$$u+��p�  u#��L$#=  �\$t=  u\��uX2���	  2�=  �L$#uց��   u΍�$�   R�D$�{A������t#h��h��h�  h���K� ��2��	  ��PS���҄�t���PU���҉D$,�\$0�\$@�\$D�\$8�\$��t$4��P����3�;L$0�	  w
;D$,�	  �T$0;�rBw;D$,v:+D$,�Q�L$8P���������  �L$4��P��3�9D$,��  9L$0��  h   ��$�   j P�,i �|$@�w��R���΃���$�   P�Oh   ���ҋ؁�   �\$`�ws�D$�D$(���D$<�;؉D$L�Y  ��   �M  �D$,���   ��$�   �T$0 3�9�$�  ��;ϋ�l$�  �׋�+Ѓ��  �|$ ��$�   t)��$�   ��$�   �L$��$�   �T$�D$�L$�'��$�   ��$�   �T$��$�   �D$�L$�T$��$�   ����  ��$�  ;L$��   �   �C�;��s  ���$    ��T$R��4�   �L$�׉l$�����L$����t"9�$�  t�D$,�C��T$0 ��;�v��!  �|$ ��������  ���  9�$�  ��  �D$ ���������|$(�\$�l$ ��u$�D$P�L$ ��$�   �����l$$�\$ �����(�L$Q�L$p��$�   ����������t
�\$l�\$3������  ���{  ���q  �T$<3ɍT�$�  �\$P�$�  �l$T;��0  r
9T$�$  �T$(�B3�;D$�*  ;��"  �l$8���  ;��L$�	  ��+ƃ���  8L$t�N�F�L$�N�D$����F�L$�N�D$�F���D$�L$��  ���9\$��  ���\$�\$ ��u�L$Q�L$ ���P����L$$�D$ ���!�T$R�L$\������������a  �D$X3Ʌ��S  ���K  ��u!�D$,ÉD$@�D$0ÉD$D�D$8   �&  �D$8   �  �|$ �\$t3�D$(h��  VPS��$�   ����������  ;���  ��+ΉL$H��$�  3Ʌ���;ǉL$��  ��+Ѓ���  �|$ t�H�P�L$�H�T$����P�L$�H�T$�P���T$�L$�l  9t$�b  �����|$(�l$�t$ S��u�L$ �	����t$$�l$ �����$�   ���������  �l$|3����  ���  ����  �|$ �l$d�t$hto�D$(�L$H���3���;D$P��  ;L$T��  �T$`�t$4j R����������  ��P����3Ƀ��;D$,��  ;L$0��  �D$�  �L$(����   �L$<3��$�  �$�  ;��V  w;��L  �T$L3���;L$T�8  r
;T$P�,  �|$' ��   ;��D$    �  ��+Ѓ��  �|$ t�H�P�L$�H�T$����P�L$�H�T$�P���T$�L$��  �|$q  ���  �|$(�t$��Vu	3��`������$�   �����������  ��t$;��D$    �j  ��+ȃ��]  �|$ t�P�H�T$�P�L$����H�T$�P�L$�H���L$�T$�  �|$� �  ����|$(�L$�L$ V��u�L$ �����T$$�t$ ������L$|�8����������  �t$x3҅���  ����  ����  �D$<�L@3��$�  �t$p�$�  �T$t;��|  w;��r  �\$(3��K���� ;D$h�U  r
;L$d�I  ��$�   R�39���T$��h�� ��$�   USR���#�������������  ;��  ��+�;��D$    ��   ��+ȃ���   �|$ t�P�H�T$�P�L$����H�T$�P�L$�H���L$�T$��   �|$�� ��   ������L$�L$ u�T$R�L$ ���7����T$$�L$ ����L$Q�L$`����������tL�L$\3҅�tB��|>��r8;�$�  r/w	;�$�  r$3�t$L�����;D$t�D���w
;t$p�8����|$ ������|$8u�D$D�L$@PQ�L$<������D$���$�   �L$43�PR������D$]��$�  _^[3��[ �Đ  �( ���������j�h{�d�    PQ�  3�P�D$d�    h(  ������D$���D$    t���{����L$d�    Y���3��L$d�    Y������������V�t$��th�W���K�����t��^�3�^����������������j�h��d�    PQSVW�  3�P�D$d�    ��h(  ������D$���D$    t����������3ۅ��D$����t'V���̷ ���   ���   ���   �   ���   �ËL$d�    Y_^[�����������V�t$��WtTh�W���z�����tD�|$��t<h�W���b�����t,V���V� ���   ���   ���   ���   �   �_�^�_2�^��������������V��������D$t	V� ������^� �̀y0 tS�A(��~L�I$��V�t���t<�~ S�\$W�|$t�VWSR��t ��f�F�~ t�FWSP�`v ���F_[^� ����VW�|$������   ��x@  u#h��hx�h(3  h���y ��_2�^� U�l$����   ��PUW��;�uUW���A���]_�^� �F   t	��u��tI�~ u'�~ u!�~ u�~ u�~( ~�~$ u	��x@  thL�hx�hf3  h���x ��]_2�^� h�hx�hm3  ��_�^� ��������������SVW�|$2ۅ�����   ��x@  ��u$hH�h,�h}3  h���(x ��_^��[� U�l$��tD��BUW��;�uUW���N���]_^�[� h��h,�h�3  h����w ��]_^��[� h��h,�h�3  ��_^�[� ������̃��  3ĉD$SUV��F�n;�W�|$,��   ���Ɂ�   v��|�nff ;�}�ȍ����   ~� �F����   ��+ȸgfff���������xi;�}e�L$�����9^��G�O�T$�W�D$�G�L$�T$�D$ }S�������F�V�����L$��T$�P�L$�H�T$�P�L$ �1;�}S�������F����F����W�P�O�H�W�P�O�H�F�L$$_^][3��V ��� �j�h�d�    P��SVW�  3�P�D$d�    �ً{��xP����+�����I �Cj<�j P��Z �K��ΉL$�L$�D$     t�2�������<���D$ ����}��C    �L$d�    Y_^[��������̃�SV��F�V;�W�|$ ��   ������   v��|� � ;�}�ȍ����   ~� �N��to��+���xf;�}b�L$�
b 9^��G�O�T$�W�D$�L$�T$}S���b?���F�L$��F_��T$�P�L$�H�T$�P�F^[��� ;�}S���%?���F���F��W�P�O�H�W_�P�F^[��� ���������V��F�V;�uE��    +���Ɂ�   v��|�Q�$ ;�}�������   ��;�}P���>����F��    +ЋFj8��j Q�Y �N�F��    +у����N��^������V��F�V;�u>��iɐ  ��   v��|�� ;�}�������   ��;�}P�������ViҐ  Vh�  j R�X �N��i��  F�����N^����V��F�V;�u;������   v��|�  ;�}�������   ��;�}P�������V��Vh�   j R�X �N����F�����N^�������������j�h�d�    PQSV�  3�P�D$d�    ��t$3�����^�^�^�^�^�^�^�F l��^$�^(�^,�\$�^0�^4�{ ��t@  �D$ ��x@  ǆ�@  �[���@  ���@  ���@  j8��<@  SQƆ|@  ��}@  ��~@  ��@  ���@  �^8�.W �����@  �ƋL$d�    Y^[��� ���������������j�hI�d�    PQSUVW�  3�P�D$d�    ��l$�E �����@  3�;��D$    t)3�;󉝔@  t���  }�ƋvP�0������;�u����5 9��@  ���@  �\$ ��[t�F;�tSP����[�^�^�^9],�u �D$ �����l�t�F;�tSP���x��^�^�^�L$d�    Y_^][�������SV��2���x@  u#h��hx�h(3  h���Hq ��^��[� W�|$��t^��PWj�҃�uWP���m���_^�[� �~ u'�~ u!�~ u�~ u�~( ~�~$ u	��x@  t-hL�hx�hf3  �h�hx�hm3  h���p ��_^��[� ���S�\$V�t$WS�6P���I�����t)��t@  u ����t��    ��Y����Q����u�_^[� ���������������������V�t$WVj���������t��t@  u
��V��N_^� ����S�\$V�t$WS��    P��������t3��t@  u*��t&�K��Y�Q��Y��Y�Q�����Q����u�_^[� ����������������������̋D$Pj����� �S�\$V�t$WS��    P���5�����tM��t@  uD��t@�K��Y�Q��Y��Y�Q���Y�Q�Q�Y�Y�Q�Q���Y�Q����u�_^[� �������������̋D$Pj�t���� ̃�S�D$Pj�D$    ������L$Q�L$�������D$�T$���[��� ����̋D$Pj�$���� �VW�|$Wj��������t��Wj�������_^� ���������̋D$Pj������ ̋D$Pj������ �VW�|$Wj���������t@�GPj��������t/�O0Qj��������t�WHRj��������t��`Wj���|���_^� ������̃�V��W�L$蠁���|$$W��������tF�ǀ   Wj���@�����t2�D$Pj���.�����t �L$Qj��������t�T$Rj���
���_^��� �̋D$Pj������ �S�\$VSj���`�����t_W�{Wj��������tL��t@  u
��W��O��t5�{Wj���������t$��t@  u
��W��O��t��Sj�������_^[� �������̃�SVW�|$ Wj��������؄��K  �GPj�ΉD$(������؄��0  �GPj�ΉD$�����؄��  �GPj�ΉD$�����؄���   �GPj�ΉD$�p����؄���   �GPj���Y����؄���   �GPj�ΉD$ �>����؄���   U�oUj���&����؄���   �?��|��<~2ۋL$$���|��<~2ۋT$���|��~2ۋD$� ��|��~2ۋL$���|��~2ۋT$���|��~2ۋE ��|=n  ~2����uh��h��h�  h���k ��]_^��[��� ������������QSVW�D$Pj���D$    �V����؄���   �|$��   th��hP�h'  �T��va�F(��~Z�N$���D���tL�@   �uC�H�ɋp|��r�Ǻ   ��;�|&;�v h �hP�h6  h����j ��2�3��D$��t�8_^��[Y� ��������{��������������SV�t$�ً��
���D$P���D$    ������tBW�|$��v8W���������q��PW��������؄ۋ�t���W����_^��[� �	����_^[� ��SUV�t$�FW3�;ǋ�t�Niɘ   QWP��N ���T$Rj�͉~������؄�t0�D$P���X��9|$~��tU��������������;|$��|�_^]��[� ���������SUV�t$�FW3�;ǋ�t�Niɐ  QWP�LN ���T$Rj�͉~�x����؄�t0�D$P������9|$~��tU���$������]> ��;|$��|�_^]��[� ���������QSUVW�|$�G3�;Ƌ�t�O��QVP��M ���T$Rj�͉w�t$ ������؄�tW�D$;�~OP���PX��9t$�t$~=��    ��t3���ud����V���K�����t��V���<����؋D$��;D$�D$|�_^]��[Y� ���������������V�t$�F��W��t�NQj P�%M ���T$Rj���F    �D$    �E�����t4�L$��~,Q���q���FP�D$P���������t�L$��|;N�N_^� ��������V�t$�F��W��t�N��Qj P�L ���T$Rj���F    �D$    �������t4�L$��~,Q���]���FP�D$P��������t�L$��|;N�N_^� ����V�t$�F��W��t�N���Qj P�L ���T$Rj���F    �D$    �?�����t4�L$��~,Q���[���FP�D$P��������t�L$��|;N�N_^� ��V�t$�F��W��t�N��Qj P�K ���T$Rj���F    �D$    �������t4�L$��~,Q�������FP�D$P��������t�L$��|;N�N_^� ����V�t$�F��W��t�N��Qj P�"K ���T$Rj���F    �D$    �B�����t7�L$��~/Q���^0���FP�D$� Q��������t�L$��|;N�N_^� ��V�t$W���N��t�F�@���Pj Q�J ���L$Qj���F    �D$    ������t7�L$��~/Q����X���FP�D$�@R��������t�L$��|;N�N_^� ������������V�t$W���N��t�F�@���Pj Q�J ���L$Qj���F    �D$    �,�����t7�L$��~/Q���T���FP�D$�@R��������t�L$��|;N�N_^� ������������SUVW�|$�G3�;Ƌ�t�O��QVP�I ���T$Rj�͉w�t$�����؄�t6�D$;�~.P������9t$~ ��t�������Pj���������;t$��|�_^]��[� ��V�t$�F��W��t�N���Qj P��H ���T$Rj���F    �D$    ������t6�L$��~.Q���Q���F�L$�PQ���������t�L$��|;N�N_^� V�t$W���N��t�F�@��Pj Q�~H ���L$Qj���F    �D$    ������t7�L$��~/Q���Q���N�D$Q�@P���w�����t�L$��|;N�N_^� �������������̃��  3ĉD$SUV�t$(�F3�;�W��t�N��QUP��G ���T$Rj�ωn�l$�	����؄�tA�D$;�~9P���#-��9l$~+��t'�D$P���m����؄�t�L$Q���=����;l$|ՋL$$_^]��[3���B ��� ����������̃��  3ĉD$SUVW�|$0�G3�;ŋ�t�O����QUP�-G ���L$�o�.����T$Rj�Ήl$�L����؄�tU�D$;�~MP������9l$~?��t;�D$P�������؄�t �L$$Qj�������؄�t�T$R���j�����;l$|��L$(_^]��[3���A ��� ����������SUV�t$W���N3�;�t�F��    +����RUQ�cF ���D$Pj�ωn�l$�����؄�tH�D$;�~@P���E{��9l$~2��t.W���������� �؄�u�F��R��P���҃�;l$|�_^]��[� ����Q�D$P�������t@V�t$��t6�L$��t)��t"h��h��h	  h���a �L$��2������^Y� ���������������������������̍D$Pj�t���� �W����t@  �uCS�\$��v5V�t$�d$ �˃���t"�VRj���:�����t
Vj���,�������u�^[_� �D$�L$�	PR������_� ���������������������̍D$Pj�t���� �W����t@  �ueS�\$��vWV�t$����˃���tD�VRj��������t,Vj��������t�F�Pj��������t�N�Qj���z�������u�^[_� �T$�D$��    RQ���U���_� �Q�$Pj�D$    �|�����t	�L$�$�Y� ����������̃��D$�$Rj�D$�D$    ��   ��� �����������̃��$Pj������t	�L$�$���� ��������������̃��D$�T$�$�$Pj�T$�c   ��� ������������̃��$Pj�B�����t�$�L$��T$�Q��� ���������{�������������̍D$Pj�d���� �W����t@  ���   S�\$����   V�t$���˃�����   �VRj���������tpVj���������tb�F�Pj���������tQ�N�Qj���������t@�V�Rj��������t/�F�Pj��������t�N�Qj��������t�V�Rj�����������g���^[_� �D$�L$��    PR���b���_� ��������������VW�|$���L$Qj�ΉD$�T�����t�W�D$Pj�ΉT$�;���_^� ������U�l$VW�D$P�}j���E     �    �+�����t$SWj�������؄�t�L$Q��$ ���E ��[_^]� ������������̍D$Pj�d���� �V��L$�$����D$�D$Pj������^� �������������̋D$Pj�$���� �VW�|$Wj���p�����t/�GPj���������t�OQj��������t��Wj������_^� ��������VW�|$�����|��<~3��D$�D$Pj�����O��|��<~3Ʉ�t�L$�L$Qj��������O��|��~3Ʉ�t�T$R�L$j��������O��|��~3Ʉ�t�D$P�L$j�������O��|��~3Ʉ�t+�L$�L$Qj���{�����t�W�D$Pj�ΉT$�b����O��|��~3Ʉ�t�L$�L$Qj���>����O��|��n  ~3Ʉ�t�T$R�L$j������_^� ��S�\$VW������������t���D$Pj�ωt$�������t��v�������PV������_^[� �������S�\$VW�����@�������v��2���w�D$Pj���D$    ����_^[� ��v&�L$Qj�ωt$�n�����t���C���PV�������_^[� ����S�\$V�s��W��}3��D$Pj�t$�.�����t��~�CPV�������_^[� ����S�\$V�s��W��}3��D$Pj�t$�������t��~�CPV�������_^[� ����S�\$V�s��W��}3��D$Pj�t$������t��~�CPV���:���_^[� ����S�\$V�s��W��}3��D$Pj�t$�n�����t��~�CP�6Q�������_^[� �S�\$V�s��W��}3��D$Pj�t$�.�����t��~�CP�vQ������_^[� �Q�D$UVW�x����}3��L$Qj�͉|$�����3���~#S3ۋ���t�T$�J�U�� ����8;�|�[_^]Y� ����������̊D$��D$�T$Rj�D$�u���� ��Q�D$P�D$ �P����L$�ɊT$tV���  �yN���F�1^�L$��t�����Y� �����������̃�$U��V�u(2����'  �M$���t����  �U �BSW���Ћ>�N3�8^�D$�\$ �|$$�L$(��  �N�ɋV(|��s"hh�hD�h
  h���X �D$,���
�L$(�|$$8^�C  8^��   �����;|$$��   ;\$(��   �T$Rj���D$ �D$ �]������D$t/f�~ �|$�\$ t h�hD�h!  �E4h���yW ���\$ �|$$�D$��v;���   r;���   h��hD�hQ  h���:W �L$8��QW���J����  �D$�8^ts�����Ã� ;|$$�D$0uU;D$(uO�F�L$Qj�͉D$��������D$�l����D$9D$�T$0�|$�T$ �N���h��hD�h9  �)����D$�4����D$�2����T$(;�r4w;�v0h@�hD�hW  h���uV �T$8��RW�������   ;�u;���   ;�u;�tw�}u�Euk�{�  �ȋE��
   ���D$��gfff����������+ʃ�	t	��	t;�)9D$#�|$8 uh��hD�hy  h���V ���D$�L$(;�rw;�v+��QW���:����;�wr;�s+��SP��衹����u�D$�M(�E �P�u ��Q���ҋF��_[~.�N���D���t �x u�x t�   �E0�D$^]��$� 3��E0�D$^]��$� �������������SUV�t$�F2ۅ���tP�������F    �V�    �    �E(����   �M$��W�|�����   �G�� t,�O������t�O�ɋG|��s3�3�QP��������G�OPQ��諵���؃���tV� tP� |J� vB�U �B����3�;u2;Ou-�O�O�M0���ٹ����V�����L$��P�AV���������_^]��[� ���W���2|�D$Pj�{���_� �D$��SVy= @�t= @�t=&  �t=q  �u6�L$�T$QR�t$�D$    �6������؋�Pj��������u<^[_� �L$�T$QR�t$�D$    谴�����؋�Pj���O�����u^[_� ^��[_� �������������QV��~2|�D$Pj����^Y� �|$ S�D$    w�D$r���w�D$��&h<�h,�h[  h���S ���D$    2ۍL$Qj��������u[^Y� ��[^Y� �����������̃��y2V�D$    �D$    |�D$Pj�����t$�T$��T$Rj�D$    �|�����t�T$3���t�L$��t��q^��� ����������QV��~2|�D$Pj����^Y� �|$ �D$    w"�D$r���w�L$Qj�ΉD$�����^Y� h<�h,�h[  h���R ���L$Qj���D$    ����^Y� ������������̃�S3ۃy2V�\$�\$|�D$Pj�����T$�ȋD$�a�D$��y= @�t= @�t=&  �t=q  �u&W�T$Rj�\$ 3�3��Z�����:�t�t$�׋�_��D$Pj�\$�9����ȋD$�:�t�t$;�t��V^��[��� �������QV�t$W�����D$    �8����D$Pj���������t9�L$��SQ��������������T$PR�������؄�t�D$P���0�����[_^Y� �������QU�l$�D$Pj���D$    ������u]YËD$��VW�x��t���W���������t*Wj V�5 �L$��VQ��������u;�t	V�����_^2�]YËT$�L$V�2 �e���;�t	V������_^�]Y��U����j�h��d�    P��`SVW�  3�P�D$pd�    ��L$<艪 ��x@  �D$x    uh��hx�h(3  �   ��P�L$Qj���҃�uB�D$Pj��������D$<t<uq��x@  �؉\$$��   h��hx�h(3  �  �~ u'�~ u!�~ u�~ u�~( ~�~$ u	��x@  thL�hx�hf3  h���'O ���L$<�D$x�����S� 3��L$pd�    Y_^[��]Ë�R�D$Pj���҃�uF�D$Pj���+����D$��t<t<u���x@  �ȉL$ ��   h��hx�h(3  �  �~ u'�~ u!�~ u�~ u�~( ~�~$ u	��x@  thL�hx�hf3  h���]N ���L$<�D$x����艩 3��L$pd�    Y_^[��]Ë�R�D$Pj���҃���   �D$Pj���]����D$<������L$��Qj�Ή|$4�������������t@  u�D$�T$�T$�D$�D$;�������D$Pj���`�����������D$��t<t<�p����L$Qj���6������L$<��   �D$x����譨 3��L$pd�    Y_^[��]Ã~ u'�~ u!�~ u�~ u�~( ~�~$ u	��x@  thL�hx�hf3  h���M ���L$<�D$x�����>� 3��L$pd�    Y_^[��]��`��PS���;�����������L$T�j`��PS���!����������j,�������D$0���D$xt�L$3�9T$ Q��W��RS�i������3ۃ��D$�D8��D$x �\$0�D$�D$ ��   ��x@  uh��hx�h(3  �a��R�D$Pj���҃�u�D$Pj���r����I�~ u'�~ u!�~ u�~ u�~( ~�~$ u	��x@  thL�hx�hf3  h����K ���L$4Qj���)�������  �C�D$4��T$��  ��   yJ���Bt!�L$,�����|���y�D$4�����X�u��D$���;��D$(%�D$4Pj���������t�K�D$4����;|$(~�;|$(�2  �|$|)�L$;�}X�S��+����    �D$4�����X�u��7;|$}1�D$4Pj���[�����t�K�D$4����;|$|��
;|$��   �|$  t�T$$���T$(��D$$�D$(�D$3���~,�W����z���L$(PQ����������D$t	��;�|��;�|x�|$  t>�D$3���~3�|$$V���z����3Ʌ�~�ȃ�;����\��|��D$�؃�;�|у|$,uC�D$��u9�C�@�����z*�[�����C���[���t��Bj�����D$0    �L$<�D$x�����%� �D$0�L$pd�    Y_^[��]���������������U����j�h��d�    P��`SVW�  3�P�D$pd�    ��3��L$<�|$ �#� ��x@  �|$xuh��hx�h(3  �   ��P�L$Qj���҃�uP�D$Pj�������D$<t<uy�ȍT$R�L$(j���������t`��x@  u}h��hx�h(3  ��   9~u"9~u9~u9~u9~(~9~$u	��x@  thL�hx�hf3  h���H ���L$<�D$x������ 3��L$pd�    Y_^[��]Ë�P�L$Qj���҃�u=�D$Pj��������D$<|��؃���x@  �\$(u}h��hx�h(3  �  9~u"9~u9~u9~u9~(~9~$u	��x@  thL�hx�hf3  h���H ���L$<�D$x�����.� 3��L$pd�    Y_^[��]Ë�R�D$Pj���҃���   �D$Pj�������D$<������L$��Qj�΃��B������������t@  u�D$�T$�T$�D$f�D$f= ��������L$Q�D�j�ΉD$<�������������   9�t@  u�D$�T$�T$�D$f�D$f;��\�����x@  ���D8��D$8u}h��hx�h(3  ��   9~u"9~u9~u9~u9~(~9~$u	��x@  thL�hx�hf3  h���F ���L$<�D$x�����ۡ 3��L$pd�    Y_^[��]Ë�R�D$PS����;�u�D$PS�������D$<uu�\$ �{�~ u'�~ u!�~ u�~ u�~( ~�~$ u	��x@  thL�hx�hf3  h���F ���L$<�D$x�����>� 3��L$pd�    Y_^[��]�<u�D$    ��x@  uh��hx�h(3  �j��R�D$PS����;�u�D$PS��������D$<uu�\$ �{�~ u'�~ u!�~ u�~ u�~( ~�~$ u	��x@  thL�hx�hf3  h���PE ���L$<�D$x�����|� 3��L$pd�    Y_^[��]�<u�D$    �L$QS���������L����D$��t<t<�8����T$RS���������#����D$��t<t<�����D$PS���l�����������D$��t<t<t<������L$QS���?�����������D$��t<t<t<������L$<�X���\$$PS��������������L$T��W��PS���������}���j@�������D$0���D$xt(�T$8�L$4R�T$,Q3�9L$(W��R��QR���\� ���3ۋC(�L$4�T$(P�D�P��Ƅ$�    �\$8�2������  �K,�T$8Q�D:�P����������   �|$  t�L$$���L$(��T$$�T$(�|$4 �D$    ~W�I 3�9|$8~/�D$WP����E �L$(PQ��������t��;|$8|��;|$8|�D$��;D$4�D$|��
�T$49T$|g�|$ us�|$4 �D$    ~d3�9t$8~6�|$$�D$VP���E ��3Ʌ�~����;��L���\��|����;t$8|΋D$��;D$4�D$|����Bj�����D$0    �L$<�D$x������ �D$0�L$pd�    Y_^[��]�����������QVW�|$�D$P��j���D$    �A�����u_3�^Y� ���   Q���������t�W���   �g!��_��^Y� ��������������V�t$V�������t&�>�   th��h��hb2  h����A ��2�^� ������̋D$VP�������L$3����@  ���@  ���@  ���@  �,����@  ��^� ���j�h؈d�    PQVW�  3�P�D$d�    ��t$�,�3�9��@  �|$t�H����@  P� �����Ή��@  ���@  ���@  ���@  �D$����������L$d�    Y_^��������j�h�d�    PQSUVW�  3�P�D$d�    ��t$j�����|$(3�;��\$ �T����@  ���@  ���@  ���@  ���@  ���@  ���@  ���@  vh�l$,;�t`8\$0t,W������;É��@  tWUP�!) �����@  ���@  ����@  9��@  t �L$4Q�Ή��@  �0����T$8RV�9 ���ƋL$d�    Y_^][��� ����������V�񋆘@  ���T�t	P��������^����������������V��F�V;�uC����+��Ɂ�   v��|�*"" ;�}�������   ��;�}P���2�������+ЋF��Q���+
���N�F����+у��N��^���̃� SU�ًC�k;�V�t$0Wul������   v��|� @ ;�}�ȍ����   ~� �K��t*��+���x!;�};�   �|$�}R���?.���t$�;�}R���-.���{��{�   �C_^][�� � ���������������j�hA�d�    P��SVW�  3�P�D$d�    ���_��x`��i��   ���    �O��V �Gh�   �j P��" �O��ΉL$�L$�D$     t� �����   ���D$ ����}��G    �L$d�    Y_^[���������SUVW�|$����}V3�9n�  �~��x%��i��   ��    �N�� �����   ;�}�N��PUQ����_�n�n�n^][� �F;�}v�N��PWQ����3�;ŉF��   �N��+�i��   i��   R�UQ��! �F��;�}*�؋�i��   +荛    �F�P��賳�����   ��u�~_^][� ~Y���;�|*��+�i��   ���荛    �N��� ���   ��u�9~~�~��F�RWP�Ή~��3�;ŉFu�n�n_^][� ������������j�hq�d�    P��SVW�  3�P�D$d�    ���_��xE�O�4�    �������G��     �OΉL$�L$�D$     t�������D$ ����y��G    �L$d�    Y_^[����SVW�|$����}@3�9^��   �~��x�F���T�����y���F�RSP����_�^�^�^^[� �F;�}Y�N��PWQ����3�;ÉF��   �N��+���R��SP�:  �^��;�}�N��R���R�����;�|�~_^[� ~J�X�;�|���$    �F��������;�}�9~~�~��F�RWP�Ή~��3�;ÉFu�^�^_^[� V�������D$t	V�k�������^� �̋D$Pj�T���� ̋D$Pj�D���� �VW�|$Wj���0�����t@�GPj��������t/�O0Qj��������t�WHRj���������t��`Wj�������_^� �������VW�|$Wj���������t��Wj������_^� ����������VW�|$W���2�����t�ǈ   Wj������_^� ��������̃� VW�|$,W���/�������   ݇�   �D$P�\$j���O�����tj����L$�$Q���� Pj���-�����tH�@+���T$�$R����� Pj��������t"��$���D$�$P����� Pj�������_^�� � ��������̋D$Pj������ �Q�D$UVW�x����}3��L$Qj�͉|$�����3���~&S3ۋ���t�T$�J�U�ͨ�����Ø   ;�|�[_^]Y� ��������Q�D$UVW�x����}3��L$Qj�͉|$����3���~#S3ۋ���t�T$�J�U轩������<;�|�[_^]Y� �����������Q�D$UVW�x����}3��L$Qj�͉|$�;���3���~#S3ۋ���t�T$�J�U�������� ;�|�[_^]Y� �����������Q�D$UVW�x����}3��L$Qj�͉|$�����3���~&S3ۋ���t�T$�J�U� �����   ;�|�[_^]Y� ��������Q�D$UVW�x����}3��L$Qj�͉|$�{���3���~&S3ۋ���t�T$�J�U� ���Ð  ;�|�[_^]Y� ��������SU�l$W����������D$Pj���B����؄�tC�L$VQ������3�9t$~%��$    ��tW���T������}�����;t$��|�^_]��[� _]��[� �SU�l$VW�}����}3��D$Pj�|$����3���~ ��$    ��t�M��P���������;�|�_^][� Q�D$SU�h3�;�W��}3�L$Qj�ωl$�Y���;�\$~^V��tX�T$�r�Vj���9�����t/�FPj��������t�NQj��������t��Vj�������L$����;͉L$|�^_][Y� �����������̋D$��SU�h3�;�W��}3�L$Qj�ωl$����;�\$~V��ty�T$�r�Vj��������tP�FPj���������t?�NQj���������t.��Vj���D�����t�T$�B�L�T$R�L$j���C����L$����;͉L$|�^_][��� ������̃�SU�l$$�EVW3�;ǋ�t�M��QWP�� ���L$�}�! �T$,Rj�Ή|$4������؄���   �D$,;��}   P������9|$,�|$~k�I ��td��D$P�\$j�Ή|$(�4�����t%�L$Qj�������L$;�u�|$ �	��u�L$ ����t�T$R��蹾���D$��;D$,�D$|�_^]��[��� �����������̀|$ �T$R��j�D$������ ����̋D$�T$Rj�D$������ ���������Q�D$S�X��U��}3ۍL$Qj�͉\$�������t4��~0V3���~(W3���t �T$�B�Pj���C������ǀ   ;�|�_^][Y� �������������̃�V��N(2�����  �V$��W�|�����  8GS�:  8Gt^�O�D$�D$�D$PjQ��. �Ѓ��D$Pj�ΉT$����f� �D$tH�F4h�h��h  h���23 ���&� t�O�T$R�L$j��������D$��D$��P���F0 �ҋ���3�;�wr;�sh��h��h)  �lU��+�ǋ�3��~2��3ɍ�   ��QP��讖����tWU���1�����u�D$WU��������u�D$ ��B����;�]t(hx�h��h@  h���`2 ���D$ ��D$�F(�V �R�~ ��P���ҋG��[~�O���D���u��B����3��F0�D$_^��Àx u�x t�   �F0�D$_^���̃�SUV��F0��D$�BW�F0 �ЍL$Q3�j�΋�3ۉ|$ �|$$�|$������t�\$���D$t�T$RS�������D$��P����3�;�rw;�v+��QP���r�����u�D$�D$�F0�D$$��t��D$(��_^][t�L$�T$��P�D$��� ������j ������������̃� �T$,3�SU�D$�D$�D$�D$�D$�D$�D$ �D$$�D$,��L$03ۅ�V�D$�L$�T$�sxJ;�u9utA�M;�u�   t�D$$f�t$&�"=�� tR=  t;;�t� �  t	�\$(�D$%�D$ �E �P����8\$$�D$�\$u*8\$%u$3��";�u��D$$f�t$&��;�u��D$$f�t$&빋�9],�E0uj�E,=�   �u }]�~�   ~�F�   �N��Ph�   Q����;ÉFt.�N���   }��   +���R���SQ� ���F�   ��^�^�D$P�M �h���^]�[�� � �������������VW�|$W��������u#h��hl�h�  h���/ ��_2�^� �N;�t#h4�hl�h�  h���[/ ��_2�^� �   9Fu-�~( ��   h��hl�h�  h���$/ ��_2�^� ��
u�~�����   ��u�~|l���   ��u�~�l���   ��u	�~6��|z��u	�~&��|l��u	�~�o�|^��u	�~���|P��u	�~\��|B9F(t#h��hl�h�  h���. ��_2�^� �N �Σ����t9xuj �������_�F    ^� hX�hl�h�  h���7. ��_2�^� �������������h  �f���������V��~uq�~t'h0�h�h�  h����- ���F    2�^Ã~( t'h��h�h�  h���- ���F    2�^Ë�Pj �҄��F    ��^�h  �����^����������̸   9At
h  ���������������̃y��h  ����������������̃y��h   �}���������������̃y��h"  �]���������������̃y|�y�o�|h#  �7���ð���̃y��h!  ����������������̃y|�y���|h%  �����ð���̃y|�y\��|h&  �����ð����h  �����������h  ����������SVWh  ���������@  ����t2Ǉ�@      3���t"��I ���  }�ƋvP�����������u�_^��[��������������V���X����D$t	V�K�������^� ��V�񋆘@  ���T�t	P���������]����D$t	V��������^� �������V��N�V;�u>��i��   =   v��|�x=
 ;�}�������   ~�	;�},P���W����"i��   N�7� �Ni��   NQ��賡���N��i��   F���N^��������������V��F�V;�uN��    ��   v��|�  ;�}�������   ��;�}5P�������N�F�����N^ËV���
����N�F��R���i����N�F�����N^���������V��~ t�j �������u�F^������VW�|$W���2�����t�ǈ   Wj������_^� ���������SU�l$W�����p����D$Pj�������؄�tC�L$VQ�������3�9t$~%��$    ��tW���D������}� ��;t$��|�^_]��[� _]��[� �SUVW�|$���������D$P3�j�͉t$�{����؄�t4�D$;�~,P���e���9t$~��t���d���P��謾����;t$��|�_^]��[� ��������Q�D$SU�h3�;�W��}3�L$Qj�ωl$�����;�\$��   V����   �T$�r�Vj���������ts�FPj��� �����tb�NQj��������tQ�VRj���n�����t@��Vj���}�����t/�FPj���������t�NQj���������t��Vj���*����L$���� ;͉L$�X���^_][Y� ������������U�������ESVW�x3�;��ى|$}�t$���L$Qj�ˉ|$�����;��t$~O��tK�U�B�0�|0��\$�D$Pj���]�����t�L$Qj�ˉ|$�����L$����;L$�L$|�_^[��]� ����������V�D$P��j�F0 �m�����t,�L$S�\$W�|$WSQ���a�����t�T$WSR���_���_[^� ��������̃�SUV��W�~�L$3�Q�ǃ�j�Ήl$�l$$�l$(�F0 �F�l$������t�T$�T$���؉~��   �|$���  ��  �D$PW�Ήl$�l$ �������S  �T$ ;��G  
9l$�;  3Ƀ~2��3�;Ѝ�   �!  w
9L$�  ��B���ЍL$Q�΋�3�������؋B����3Ʌ�w��vN;�rJw;�vD+��QP���o�����u32�3�D$(;�t�L$��D$,;�t�T$�L$ ��H_^]��[��� ��tˋ|$ �l$WU��裉����t[��B����3Ƀ~��B���Є�u2�D$�  �(;D$u;L$th��h��h�  h����% ��WU���Ɖ���؄��S����L$ �T$�D$QRP���������6���h��h��h�  h���% ��2ۉl$�����L$QW�������؄�������T$ �D$RPW���/�����������������̃�SV��L$3�2�;�u&h|�hX�h�  h���% ��^��[��� ��y&h�hX�h�  h����$ ��^��[��� W�|$;�u'h��hX�h�  h���$ ��_^��[��� U�l$$;�u(h��hX�h�  h���$ ��]_^��[��� ��E �D$ �D$�D$�D$P�L$$Q���j����T$;T$ t*hP�hX�h�  h���7$ ��]_2�^��[��� 3�9D$3|�|$s*h�hX�h�  h����# ��]_2�^��[��� �D$ �D$�D$�D$P�L$$Q���^����؄���   �T$;T$ u]�|$ |V�|$rMWj��耳���؄�t[�?}h��hX�h�  �6Uj���Z����؄�t5�}  }8h��hX�h�  �h0�hX�h�  h���D# ��2�j ������]_^��[��� ���������́�D  �  3ĉ�$@  SU��$T  V��$T  3�;�W��u�s2�r��|
��2}�4����2~h��hT�h�  ���|
��|>��2}>h(�hT�h�  h���" ��2���$P  _^][3�� ��D  � ��2|�gfff������������+�u��_4�_蔴  j@�T$SR�G�w�� ����}�2   V�D$h�P�� ���L$Qj ��賩���؄��C  j j j���<����؄��,  ��t$�}  t�ōP�I �����u�+�UP���l����؄���   h   �T$Tj R�Q ��  P�D$`h��P�f �D$h��������H����u������������Pf����H���f�P�H�D$P�����H����u������������H�P�D$P�����I �H����u�f�K�Kf��P�D$P�P�����u�+��DP���LP�L$PQ��P���u����؋�������u2ۊ��$�����������������̃�D�  3ĉD$@�T$HSUV��L$XW3����3�;׉T$�L$(�}4�}�}�|$�D$�D$ �t$$t�:�1���3�2���x@  �D$,�D$0�D$4�D$8�D$<�D$@�D$D�D$H�D$Luh��hx�h(3  �^�E �P�L$,Qj ���҃� u�D$,Pj ���K�����C9}u"9}u9}u9}u9}(~9}$u	��x@  thL�hx�hf3  h��� ���ۈ\$��  j�L$0h��Q��% ������   �D$ 3���I ��x@  �   �t$-�|$,�tP�U �R�D$KPj���҃�u[�D$KPj��蔥��j�L$0h��Q�_% ��������   ��   r��	  h��hx�h(3  h���� ����  �} u+�} u%�} u�} u�}( ~�}$ u��x@  ��  hL�hx�hf3  h��� ���  �t$$�]�D$3��   ���|, uN���� |�|$ �g  �D$;ǉut�0�T$R�D$P����������D$�%  �|$t_�D$ �  �� }��T$K���|$ �  ��u��Xu�2�T$K�L,��0|��9�Ƀ��� �4��tq�|��o����D$ ��  �D$ ;���   �t$;���   ;�|-����� v#h`�h8�hH  h��� ���D$ �t�\$(�NQ�ˋ�芞��V������V���:������  �@���PV��������~2���V�������8 tV�������8uV��������������  �W��艥��3�W���������'����|$ ��   �}��   �U �B���Ћ�3��d$ �L$Q�T$R�����������   �D$=  w-=  ��   �ȁ�   ��   ��   ��   ���   =  ��   =  ��   =  r=  ��   %  ��=   u3h��h8�h�  h���" ��9|$�E   t
�T$�   �}u#�E �P����3�;�rw;�v+��QP�������L$P�D$_^][3���� ��D� =% @��t����D$P�L$Q���j�����t�W���N���������������j�h��d�    P��$SUVW�  3�P�D$8d�    ��|$H���E    � �E �P���҃}���t$,�D$ �D$ �D$ �D$ �D$ ��   �D$0P�L$$Q���D$(    ������؄���  �|$   uU���= ������D$j ��������u2��D$�|$   ��  ����  �T$0R�D$$P���D$(    �^����؄�u��~  �U �Bj ���ЍL$03�Q�T$$R�͉D$(�D$8�D$<�(����؄��8  3��D$ =  ��  �Q  ���  - @ ��  -�����  �GXPj���D$!�&����؄���  �O`Qj�������؄��t  �WdRj��������؄��]  �GhPj�������؄��F  �OlQj���ʩ���؄��/  �T$$Rj��販���؄��  �D$$;��  ��P�3������D$(��Pj V�A� �L$4��VQ���A����؄�t	V�OT����V�<������D$$    �  �D$4���t$0��  ��@B v!h$ h  hG  h���9 ���  ���x  	���m  �L$���S����VR�L$ �D$D    �����V�L$ �T���V�L$ 誠���L$�  计��PV��腟����~8���V�L$ 脠���8 tV�L$ �u����8uV�L$ �f����������  �W�L$ �����L$�V��������<  �> t=��$    j
h��V� 0 ����t
���> u���F
��
��t< 
�F����u�3�8��   �<0(t���<0 u��'���0 ~��$    �0�� ~��-u�0 �����> ��   j
h��V3��/ ����uk�L$Hh�����   ������F
���~
t< 
�G����u�<0|<9~<.u������t&< "� �G����t�I < ~<-u
�G����u�> t�L$HV���   艿����t�? t�L$HW���   �p����L$�D$@����������|$H�u  �D$ Pj���D$ �t$(�����؄�te�D$ ;�~L��P�x����L$$��Q��j V�� �T$0��VR��膝���؄�tV�������V�������D$     3���t�GP��薩���؄ۉt$(��   �L$(Qj���j����؄���   �T$ Rj���R����؄���   �D$ ;�~K��P��������D$$��Pj V��� �L$0��VQ�������؄�t	V�O�V���V��������D$     ��t`�W,R��������؄�tO�D$(Pj���ҥ���؄�t;�OPQj��迥�����*=  t=% @�u�D$��Wp�B$�OpU�Ѕ��È\$3�V���'�����u2ۀ|$ t�|$ t�|$ uC�|$ u<��t8�L$0Q�T$$R�͉t$(�t$8�t$<������؄�������t$,���|$ tL��t$,�E �P����3�3�;�u;�t0;�rw;�v+��QP���y���;�wr;�s+��RV���x���ËL$8d�    Y_^][��0� ������̃�V��~u�L$V�za��^��� U�l$SW�D$P�L$ Q���D$$    �3����؄�t/�|$��  u
V���9a����j ���������t��  t��u�_��[]^��� _[]2�^��� ������j�hӉd�    P��SUVW�  3�P�D$,d�    ��L$�^����D$$P�L$3�Q�͉|$<�D$ �|$ �������\$<tr� @ �9t$t'W���b�����tZ�T$$R�D$P�͉|$ �Y�����u��?jp�������D$<;��D$4t	���%����3���E�H�M�P�D$8 �i  �D$9;��  �T$$R�D$P���D$ �|$ �|$,�|$0��������N  ���t$�� @ ��   �� @�th��3 @���   �D$$���L$(u;�t6��u;�t�j������W�A����   �j������j�*����   �W������W�����   �L$$Q�L$$������R�����u�D$<Pj�͉|$D脢���D$<='  w<P�L$ �����L$�V���P�L$ �̎��P���$�����t/�L$�g����P������hd h@ h7  h���D ��W��蹹����t1���t'�L$$Q�T$R�͉|$ �|$,�|$0�������������D$W���|�����u�D$��|$ u�;���   ��Pj�҉;�   9;��   ��x@  ��   9}��   �}��   �L$������L$���e�������t$��� ��|]�G�=�   wS��tO�> tJ�OQj�������V�V����Ė �N��D$WPQ�~��� �V� ���@  �F�����@  �L$�D$4���������D$�L$,d�    Y_^][��$� ������������j�h �d�    P��TSUVW�  3�P�D$hd�    ����$�   3�;�t��L$8�\$軙����$�   �l$x;��O�L$<�D$����t���4���t$|;�tL�������h�   h�   h�   �N(����h�   h�   h�   �N0�כ��SSS�N$�̛���
��$    �I ��$�   ��T$<�Wt0�D$HP�L$$Q�ω\$(��������  ��$�   9T$ ��  3ۍD$HP�L$$Q�ω\$(�\$P�\$T�b�������  �D$ ;�$�   �c  =  @��  ��  = @ �  ��   =�� tw= @ ��  �L$$輋���T$$�   R�ω\$t�7����L$$讋����~+�D$|��t�Hd�:������D$$P�N�[����^$��$�   ��L$$�D$p���������  ����  �UR���v����  �|$| ��  �L$(�-����D$(�   P�ω\$t訽���L$(������t+�L$|��d诟���L$(��Q�N�к����$�   �^$�   �L$(�D$p�����_����  = @ t`=  ��  ����  �L$,觊���D$,P���D$t    �#����L$,蚊����~�L$,Q�M�Y����L$,�D$p����������  �L$0�Z����T$@Rj���D$x   �����|$@u;�D$0P��������L$0�8�����~"�D$|��t�L$0Q�H������$�   �   �L$0�D$p����聍���;  ���3  �L$D�ۉ���L$�D$p   �ʉ���D$4P3�j���D$x�\$<��$�   �J����L$xQj���<����T$4R�L$讕���L$����P�D$8P�������L$�/���Ph� �ĝ  ����up�D$x;���  ��P��������L$|����T$xVR��蝓������   �|$���   V����x��;ÉD$��   S�͉E �k��V�u������  �L$褉��Ph� �9�  ����u}�D$x;��i  ��P�������� �D$|��� �L$xVQ��������t9�|$�u*V���Mx��;ÉD$|"j�͉E ���V��������  �D$����V���������   �L$����Ph� 衜  ����ug�|$xu`�L$P����T$PRj���<�������   ��$�   ;���   �L$P�T$T�H�L$X�P�T$\�H�L$`�P�T$d�H�    �P�v�L$芈��Ph� ��  ����uW�D$x;�~S��P�������� �D$|��� �L$xVQ���������t��$�   ;�tV�H�    �,���V���������O�L$�D$p�ߊ���L$D�D$p�����Ί���  = @��  ��   = @�t^= @��  �L$H�D$L���������O  r���   �A  �L$|��t�l$H���5x4�$�E\����$�   �   �  �\$H����� u�|$L ��   �t$|��tW�D$J��PQ�Ӂ��   R�L$D�ؕ���D$8P���L\���[�����ۉ\$ �D$ }�h+�5�'�������$�}[����$�   �   �   ����   �T$J�D$H��RQ%�   P�MP�g����d=" @�t8=  �t�O�P��tL�D$���t9E t>�|$L w7�D$Hr=���w*�E �%�T$H�D$L�ʃ�������wr�����w��t�Ulj ��������t3��-����D$�j ���Ͱ���D$�T$<��$�   �W�8 t��t�O�M(�L$|��t	�WR�K[���G�D$�L$hd�    Y_^][��`� �������������j�hi�d�    PQSUVW�  3�P�D$d�    ��t$�|$(W軄���D��G�F�O�N�W�V�G�F�O�W�N3�R�N�l$$�����G P�N �D$$�����O$�N$�W(�V(�G,�F,�O0�N0�W4�V4�G8�F8�G@�^@�^d�GH�D$ �^H�GP�^P�GX�^X�O`�N`�Wa�Vaf�Gbf�Fb�OdQ������k�k�k�r����0��Nt�WtR�D$$����i�i�i������   ���   ���   �P���   �H���   �P���   �ƋL$d�    Y_^][��� ������U����j�h��d�    P��  �  3ĉ�$p  SVW�  3�P��$�  d�    �E��M�L$(��$�   �D$����3�9~(��$�  t:hh� h5&  h��� ����$�   Ǆ$�  �����s���3���  �T$R�D$P�Ή|$�g�������  � � 9\$t+j ���;������q  �L$Q�T$R���2�����u��W  ��$�   �-���L$|�$���L$4�����$�   Pj���ʖ�������  �L$|Qj��豖��������  �T$4Rj��蘖��������  �D$,Pj������������  �L$Qj���f���������  ��$�   Rj���J���������  �|$ ��  �D$4P��$�   Q�T$TR��"���D$(����$�   P��$�   Q�T$TR����$�   �$P�������������L$dQ�L$P������D$��������Au���L$l�$������h�   訩�����D$��Ƅ$�  t���N@�����3�j	��Ƅ$�   �'E����$�   R����F���D$dP����F���� �����$�E�����D$,������Au%�D$��������Au���d �����$��D������؅ۋL$�tV�\$(j j��T$R��$�   PS���D$(    ������t�C(�����|$ t�L$Q��$�   �OV����D$�R��E��j ���ȫ����u3���$�   Ǆ$�  ����諓���ǋ�$�  d�    Y_^[��$p  3��� ��]� ���j�h�d�    P��dSUVW�  3�P�D$xd�    ���G(3�;É\$ ~4�O$���l�;�l$t"�}  u9]u9]u��B���ЉD$ ��\$��L$(�\$�#���L$X�p���L$(Qj�ω�$�   �œ��:ÈD$�~  ��$�   �T$XRj��D$$PSQ���M����D$�D$X����   ��tGj 耧������$�   ;�Ƅ$�   t�T$(R���>v����$�   ��  ��$�   3���  j(�9�������$�   ;�Ƅ$�   t���,� ���3��T$(�V�D$,�F�L$0�N�T$4�V�D$8�F�L$<�T$\�N�n R�͈�$�   薮����������th0g��菪����$�   �l$�0��   �L$`�����;����A��   j8茦������$�   ;�Ƅ$�   t����� ���3��L$(�N�T$,�V�D$0�F�L$4�N�T$8�V�D$<�L$`Q�T$DR�L$0��$�   �F�5����N �P�V$�H�N(�P�V,�H�N0�P��$�   �V4�0�=j ��������$�   ;�Ƅ$�   t�L$(Q���t���3���$�   ���$�   8\$ty3�;�w9\$ vm;�ti�G(;�~�O$���D��3�;�uP�}  uG9]uB9]u=��B����3�;�r.w;D$ v&+D$ ΋��փ�������;�wr�����w�u�M�L$\Ǆ$�   ����藀���D$�L$xd�    Y_^][��p� �������������U����j�h�d�    P���  �  3ĉ�$�  SVW�  3�P��$�  d�    �E���M��$�   �L$�D$42��     �|����E������Ǆ$�      �{  �$�l�	�T$HRj�������؄��  �D$H��t	���%  �D$ Pj��������؄���  h�   �-������D$��Ƅ$�  t	���c� �3�j�ȉD$ Ƅ$�   �
� �L$L�!�  �L$LQj��Ƅ$�  �ۏ������  �T$dRj���ŏ������  �D$|Pj��诏�����{  �t$L�Nl����Q�L$ ��� �T$RW��$T  �`��������I  �L$������t$P����� �D$Pj���Ҏ��2�:�u��$�  �  �L$8Qj��貎��:�t�T$RW��$T  �����������  Q�D$�̉d$ P�0������9c���L$Q�   S���g�������  �T$�D$<PS�ω��   �Ȏ������  �D$<ݞ�   9\$Hu*�L$<QS��裎�����o  �T$<RS��莎�����Z  ����� ���h���;�Ƅ$�   }.�D$4�L$L�     �9Y �L$Ǆ$�  �����E������O  �L$4�1� 	  �T$ Rj��襍�����  �|$ u��D$ Pj��舍������  h�   ��������D$��Ƅ$�  t����� ���3�j��Ƅ$�   ��� �L$L���  �L$LQj��Ƅ$�  覍�����r  �T$dRj��萍�����\  �D$|Pj���z������F  �t$L�j����Q���� �T$Rj���ь�����  �D$8Pj��軌�����  �L$DQj��襌������   �L$D��}K��Ƅ$�   ��W �L$Ǆ$�  �����������$�  d�    Y_^[��$�  3��i� ��]� 3��D$$lI�D$(�D$,�D$0;�Ƅ$�  �D$~G�I ��$�   Rj��菌����tN��$�   P��$  ����P�L$(��/���D$��;D$D�D$|��L$$Q���� �T$4�Ƅ$�  ��  Ƅ$�  �L$$����Ƅ$�   �L$L��V �L$Ǆ$�  ��������2������D$ Pj���r�����tӃ|$ ������L$ Qj���U�����t�h�   �ǟ�����D$��Ƅ$�  t����� �؉D$�3ۉ\$�D$ �����Ƅ$�   w����	�$���	j�j���� �L$L��  �D$LPj��Ƅ$�  �Q����������L$dQj���;����������T$|Rj���%�����������t$L��g����P���:� 3��D$$lI�D$(�D$,�D$0Ƅ$�  �D$���    ��$�   Qj���ϊ������   ��$�   R��$   ���P�L$(�9.���D$�����D$|��t$�D$$P����� �L$QW��$T  �W���������   �L$����P����� �T$RW�0�������tj�L$�Ц��P����� �D$Pj��誉����tG�L$Q���� �T$Rj��茉����t)�D$8Pj���z�����Ƅ$�  ������L$4�1�  Ƅ$�  �����T$ Rj���D�����������|$ �X����D$ Pj���#����������h�   葝�����D$��Ƅ$�  	t���� �؉D$�3ۉ\$j��Ƅ$�   �h� �L$L��  �L$LQj��Ƅ$�  
�9����������T$dRj���#�����������D$|Pj��������������t$L�e����Q���"� �T$<Rj��������������D$<�D$<Pݛ�   j���Ĉ����������D$<��$,  Qݛ�   j��衈�����m���3��D$$lI�D$(�D$,�D$0Ƅ$�  �D$��$    ��$�   Rj���_�������   ��$�   P��$�   ���P�L$(��+���D$�����D$|��t$�L$$Q���i� �T$RW��$T  ����������   �L$胤��P���[� �D$PW���������tn�L$�`���P���X� �L$Qj���:�����tK�T$R���J� �D$Pj��������t-�L$8Qj���
�����Ƅ$�  
�L$$�E����T$4�2�)  Ƅ$�  
�)����D$ Pj���І�����-����|$ ������L$ Qj��识��������h�   �������D$��Ƅ$�  t���c� �؉D$�3ۉ\$�D$ ��Ƅ$�   t	��uj�j����� �L$L���  �T$LRj��Ƅ$�  賆���������D$dPj��蝆�����i����L$|Qj��臆�����S����t$L�&c����R���� 3��D$$lI�D$(�D$,�D$0Ƅ$�  �D$��$�   Pj���9������.  ��$�   Q��$   �m	��P�L$(�)���D$�����D$|��t$�T$$R���C� �D$PW��$T  �����������   �L$�]���P���5� �L$QW蚤��������   �L$�6���P���.� �T$Rj����������   �D$P���� �L$Qj��������tg�T$8Rj���܄����Ƅ$�  �����D$4�0�L$$������Ƅ$�   �L$L�
P ��$�   j j��L$$Qj R���D$0    ��������Ƅ$�  ��������	-�	`�	��	�	�	�	    ���������������j�h3�d�    P��   �  3ĉ�$�   SUVW�  3�P��$�   d�    ��$�   ����$�   ��$�   �D$0R�D$(�L$P3�P���D$ �t$,�~������n  �|$$  �  �L$P�t$�t$ �t$,�t$$�_N �L$Qj�ω�$�   芃����u�L$PǄ$�   ������N ��  9t$~�T$ Rj���Y�����t�9t$ ~ɍD$,Pj���A�����t��L$$Qj���/�����t��T$PRj��蝃����t��D$hPj��苃����t�h�  �}�������$�   ;�Ƅ$�   t%9t$$��9t$,��Q�L$ R�T$(QR����V�����3ۍ�$�   P�L$TƄ$�    �\$,蓊 ݄$�   �X�L$4�����\$D݄$�   ��ݜ$�   ܼ$�   ݜ$�   �'���D$3�;���   ��$�   Qj�Ͼ   �y������   ��t@  u��$�   ��P����H����u���$�   ��$�   ��$�   �D$�D$4�D$�L$P�K�L$H�D$T�\$8�D$�T$܌$�   �D$\�\$<�D$܌$�   �D$d�\$@� (���D$��;��H�����D$9C��  =��  ��   3�9l$ ��   ��$�   Qj�Ͼ   �5x������   ��t@  u��$�   ��P����H����u�K�(����$�   ���$�   �P��$�   �H��$�   ���P;l$ |��I3�9t$ ~A�I �D$4Pj��������t,�K�&(���L$4��T$8�P�L$<�H�T$@���P;t$ |D$ 9C ��  �|$, �#  �L$4�Q��3�9t$�  ��I ��x@  ��   ��R�D$Pj���҃���   �D$Pj���v���L$��$�   �T$ۄ$�   �P��$�   ���D$�L$4Q�K(���\$8ۄ$�   ��$�   ���\$<ۄ$�   ���\$@�<&����;t$�_����Zh��hx�h(3  �<� u'� u!� u� u�( ~�$ u	��x@  thL�hx�hf3  h����  ���C0;C��   �|$$ ��   �L$D�#��3�9l$��   ��$    �T$Rj�Ͼ   �v����tx��t@  u�D$��P����H����u��D$��$�   �L$ۄ$�   �X��$�   ���T$DR���   ���\$Hۄ$�   ���\$L��#����;l$�q������   ;Cu�D$�L$PǄ$�   ������I �t$(j ���0�����t^�|$ tW��tb�D$0�T$Lj j��L$8Qj R�ω0�D$D    �����D$��$�   d�    Y_^][��$�   3��Q� �Ĭ   � ��t��Bj�����D$ ��������̃�S3�2ۅ����L$Q�T$R�ΉD$������t(9|$t)j ���{�����t�D$P�L$Q���v�����u؊�[��ð[�������VW��	 �    ��������u_3�^Ë�艝��j �Ή������u3��; u3���_^�������������VW��  �    �<�������t>� �+�������t��荣��j �Ή�����u3�j ��賔����u3����u���t��Pj���    ��_^��������������U����j�h��d�    P��   SVW�  3�P��$�   d�    3ۍL$T�\$<�\$4�[G �}��x@  ��$�   uh��hx�h(3  �[��P�L$/Qj���҃�u�D$/Pj����r���C9_u"9_u9_u9_u9_(~9_$u	��x@  thL�hx�hf3  h���2�  ���D$/<t<��  ��x@  ��uh��hx�h(3  �[��R�D$/Pj���҃�u�D$/Pj���/r���C9_u"9_u9_u9_u9_(~9_$u	��x@  thL�hx�hf3  h����  ���D$/<�t��t<t<�I  �L$0Qj���$r����t��t@  u�D$0�T$1�T$0�D$1f�|$0�  �L$T�����PV���{���L$l�����PV���{���\$0�ۉ\$H�D$8    ��  3��D$@�D$L�D$P�D$LP�L$DQ3��ωt$L�y������q  �|$@	  u!9t$P|9t$Lv�\$D��������t$D�\$Hj ���-������&  ���-  �|$8 u2j(�������D$D��Ƅ$�   t
S����� �3�Ƅ$�    �D$4���m� ����   ���M������   ���������   jP莎�����D$D��Ƅ$�   t���% ���3ۋF�@���\$�K8� Ƅ$�    �$�<���SRj ���,���C Pj���r,���N�KH��Bj���ЋL$4S��$ �\$H��������u���n���L$4V�$ �D$8��;ÉD$8�s������t��Bj���Ћt$4��t/���a��;Ë�u�V����uFj ����� �D$<�΋�Bj�ЍL$TǄ$�   �����eD �D$<��$�   d�    Y_^[��]Ét$<������̃�,S3�UV�t$<�D$�D$�D$<��P���nw���D$<���  �yM���E�ȃ��L$$�L$Q��j�ΉD$(�x����u^]2�[��,� �T$Rj���ox����t�D$Pj���]x����tэL$0Qj����x����t��T$(Rj���x����t�W�  ��������   � ������tV�.�����j �΋�蠏����|$j ��葏����trW���������D$|W����   �  ������tL� ������tV�������j �΋��E�����|$j ���6�����tW���:�����}��Pj����_^]2�[��,� P������L$�T$HQ3�9L$R��QP���O����T$HP3�9D$R����P�Q���x8��|y�D$,��i��   sdݞ�   �D$4ݞ�   �L$�T$ QR���;5���|$$ t��_�FP   ^]��[��,� �|$( t��_�FP   ^]��[��,� ��������nP��_^]��[��,� �����UV�t$W�  ���}�����u_^]� S� �h����؄�t#�D$�L$PQV������j �Ί��������u2�j ��������u2ۊ�[_^]� ������̃�(UV�t$4W�D$P��j��3��v����u_^2�]��(� �|$|�L$Qj����u����t܋T$����wЍD$Pj���Rv����t��D$���t��t
��u�x��   ��   �t$<SVW�����3�9\$��~�I �L$<WVQ���������t��;\$|�[_^�]��(� [_^2�]��(� �������������UV�t$W�  ���-�����u_^]� S� �����؄�t�D$PV�������j �Ί�誌����u2�j ��蛌����u2ۊ�[_^]� ������������j�h��d�    P��TSUVW�  3�P�D$hd�    ��3ۍL$0�\$$�(�  �L$8�\$p�\$�\$(�\$�\$�K? �Gh�l$x�L$Qj���D$x�D$4�mt��:���  �|$�~  �T$(Rj���Lt��:��h  �D$Pj���6t��:��R  �D$�ȁ�  �yI���A�+L$x���L$8�D$�����Pj���{t�����  �L$P����Pj���`t������  �L$Qj����s��:���  �D$;�~� R�L$4蝁  �D$ �D$��\$ ;�~�L$ QP����r��:���  �\$$��������u
�D$p �  �D$$��t�P��荜��P���%���|$ ���V0�D$�^P���Y���|$x �D$$����u�L$$Q���i���D$x3�;\$}VU�����������D$xu�D$����   �wh��    R�L$4�̀  �T$,3�;֋؋�})i��   ;L$}!�od�|*Pu���������   ;�|�;L$��   �T$3����   �D$ �hf��|q��;�}j�����wd�D$,i��   �T0@�L$$i��   ����t1@u��|�Od�t@k�h�GT�T$,R�LH����u��|�Gd�T@k�h�GT�L$$Q�LH� h���T$��;��s����L$8�D$p �S= �L$0�D$p�����2�  �D$x� �\$p�L$8�/= �L$0�D$p������  2��L$hd�    Y_^][��`� ������j�h��d�    P��\SUVW�  3�P�D$pd�    �ٍL$0��~  3�L$@�l$x�l$,�l$$�l$�< �{h��$�   �D$,Pj��Ƅ$�   �|$0�/q���L$$Qj���!q���T$@Rj���q���D$XPj���q���L$Qj����p���D$;�~� R�L$4��~  �D$ �D$��l$ ;�~�L$ QP���3p��Ƅ$�   �l$�T$;T$$��   �D$8P�L$Q��Ƅ$�    �l$ �<�����t7���    �|$  �b  U���
�����t�T$8R�D$P��������uъ�$�   ����$�   tR� �%�������$�   t#V���B���j �Έ�$�   貇����u��$�   j ��螇���|$(3��u��$�   �D$��$�    �#����D$;���   �sh��    Q�L$4�}  3�;����},i��   ��;L$}"�{d�|Pu�D� �������   ;�|�;L$��   �T$3�����   �D$ �xf��|z��;�}s�D� �L� �sd�D$(i��   �T0@�L$i��   ����t1@u#��|�Kd�t@k�h�CT�T$(R�LH�&��������u��|�Cd�T@k�h�CT�L$Q�LH��d���T$��;��j����L$@�D$x �(: �L$0�D$x�����~  ��$�   �L$pd�    Y_^][��h� ���������̃�VW3�Wh �D$P��L$(WQ�Ή|$�|$ �����T$R�D$P��������u
_2�^��� �|$ uV�X�������j ���ʅ����tԋL$�9_^��� ��������j�h�d�    PQSVW�  3�P�D$d�    ��L$(j h �D$Pj Q���D$$    �������u2��L$d�    Y_^[��� � ������t�h�   �������D$(���D$    t���������3�V���D$ ��������j �Ί��������u2����u��t(��Bj��������FH����������8p���L$$�9�ËL$d�    Y_^[��� �����������j�hK�d�    PQSVW�  3�P�D$d�    ��L$(j h �D$Pj Q���D$$    �������u2��L$d�    Y_^[��� � ������t�h�   �������D$(���D$    t���������3�V���D$ ��������j �Ί�������u2����u��t(��Bj��������6G����������(o���L$$�9�ËL$d�    Y_^[��� �����������j�h{�d�    P��(SUW�  3�P�D$8d�    �D$0P�L$3�Q��3��\$0�\$�]�����u3��L$8d�    Y_][��4Á|$�� �Z  �T$$R�   U���tk�����@  �D$$%������d�D$$t	��e�%  �D$PU���Dk��9l$�  �L$ QU���-k��9l$ ��   �T$RU���k���|$��   �D$PU����j���L$;L$��   �T$,RU����j��9\$,��   j,�R�����D$;É\$@t�L$�T$Q�L$$R�T$$QR���V�����3�E�L$�T$P�D
�P���D$H�����l$��j����tJ9\$ �\$t��3�9|$~+��I W���
��PS����j����t��;|$|��;|$|�D$(   3ۋ|$S���ā����t9\$(u;�t��Bj���Љ\$���ǋL$8d�    Y_][��4�j�h��d�    P��0SUV�  3�P�D$@d�    �D$$P�L$Q3ۋ��D$ �\$�^�����u3��L$@d�    Y^][��<Á|$�� ��  �T$ R�   U���ui������  �D$ %������d�D$ t	��e��  �D$PU���Ei��9l$��  �L$QU���.i��9l$�|  �T$8RU���i���   9t$8�`  �D$<PU����h��9t$<�I  �L$0QU����h���T$0;T$8�.  �D$4PU����h���L$4;L$<�  �T$,RU���h��3�9l$,��   j@�}�����D$$;ŉl$Ht)�L$4�T$0Q�L$@R�T$@Q�L$(R�T$(QR����' ���3ۋC(�L$8�T$0P�D
�P���D$P�����\$�h������   �K,�T$<�D$4Q�L�Q���h����tm9l$t�T$���T$$��D$�D$$�|$0 ~F�D$43���~+VU����  �L$$PQ���Wh�����D$4t	��;�|��;�|��;l$0|��;l$0|�D$�\$j ���?����t�|$ u��t��Bj�����D$    �\$�ËL$@d�    Y^][��<�����QSV��2��D$    �\�����t"�L$j h�� �T$R��D$ j P�γ�V���^��[Y� ��������������j�hۍd�    P��SUVW�  3�P�D$,d�    ��D$3�Pj3ۉ|$$3�|$�|$ ��f����u3��L$,d�    Y_^][��$ËD$��|���|$ ��   �L$$Q�T$R���9�������   �|$  u������j ���~����tk��tg��u���J��u;j(��z�����D$3�;ǉ|$4t	���c� ��S���D$8�����|$ �] �ߋ|$ �L$U�M ��3�;|$�|$ �`����';|$}!��t�E �Pj���҅�t��Pj����3ۋËL$,d�    Y_^][��$������������j�h,�d�    P��   SUVW�  3�P��$�   d�    ����$�   �   ��I ���)�������y�3��D$@�D$�D$8�D$�D$$P�L$ Q��������u2���  �|$�� �s  �T$<Rj���D$D�����e�����U  �D$<��dt��eu�h�   �oy�����D$8��Ǆ$�       t	���2
���3��D$ �D$8�D$Pj��Ǆ$�   �����d������  �D$����  �l$ ��P����� 3�9t$~1����i������D$t�L$Q���~����;t$|��
;t$��  �T$Rj���Bd������  �D$���{  �l$ �� P���^� 3�9t$~6��    ����������D$t�D$P���}����;t$|��
;t$�.  �L$Qj����c�����  �D$���  �\$ ��0P����� 3�9l$~h��    �T$$R�D$ 3�P�ωt$$�9�����t=�|$	  u������j ���{����t��t�L$Q�ˉt$ ��|����;l$|��
;l$��  �T$R�   U���,c���D$�L$ P��@���3�9\$~b�I �L$ �w
�����F(PU����b����t:�NQj���hc����t)�V,R����j����t��@VU���Ic����t
�;\$|��
;\$��  �D$PU���b���L$Q�L$$��P�����3�9\$��   ��$    �L$$������L$ j���$�   �
�����F8PU���Wb������   �F<PU���Cb������   �T$$Rj���b����ty�L$$�T$(���ĉ�L$<�P�T$@�H�ΉP�) �F@Pj����a����tA�FHP����i����t2��XVU���Vb����Ǆ$�   �����L$$t"�- �;\$�2�����L$$Ǆ$�   ������, ;\$��  �L$QU���a���T$�L$ R��`������|$ �D$    ��  �\$ j����t8�����F8PU���Fa������  �F<PU���2a������  �L$$�����D$$Pj��Ǆ$�      �a�����p  �L$$�T$(���ĉ�L$<�P�T$@�Hj �ΉP�C �F@PU����`�����3  �FDPj���`�����  �FL�L$4QU�ωD$<�`�����  �|$4 �D$4P��U�ψVL�y`������   �D$4�����w%�$���	�nP��FP   ��FP   ��FP   �L$4QU���3`������   �FXPU���`������   ��`Vj���`����tv��$�   Rj���u`����ta��$�   Pj���``����tL�L$|QU���O`����t;�T$DRU���>`����Ǆ$�   �����L$$t*�+ �D$�;D$�D$�5����"�L$$Ǆ$�   ������* �D$;D$��  �L$QU���a_���T$�L$ R��p�����3�9\$��   �d$ �L$ j �������FPU���'_����t_�FP���g����tP�L$4QU���_����t?�D$4+�t+�t+�u�F$   ��F$   ��n$�F(PU����^����t
�;\$|��
;\$�  �T$RU���^���D$�L$ P���   �I���3�9\$~q��L$ j��U	�����FPU���w^����tM�NQ���hf����t>�F,PU���X^����t.�V0�D$PU�ωT$$�?^����t�|$ ��݈N0;\$|��;\$|n�L$L��( �T$LRj��Ǆ$�      �~^����u�L$LǄ$�   �����F) �2�D$dPj���V^����Ǆ$�   �����L$Lu�) �
�) �D$j ���Iu����t\�|$ tU�t$8��t^���	����$�   ��$�   j �1h�� �L$HQj R��虼���D$��$�   d�    Y_^][�Ĭ   � �L$8��t	��Bj���D$ �Ȑ��	��	��	��	��SUVW���D$P�L$Q3��ωt$谥�����  �\$$�l$ �D$=	  �  ��   =  ��   t`-  t1����  �D$(    ��  SU�����������������  �D$(    �q  SU�����������������\  �D$(    �I  SU������������������4  =  �)  �D$(    �  SU������������������  �D$(    ��   �D$$    ������t#j h�� �T$,Rj S�ωE �����   �   ����   =  w{tX=  t0=  ��   �D$(   ��   SU�����������������w�D$(    thSU������������������V�D$(    tGSU�����������������5=   r.=   w'�D$(   tSUP������������������   j ���r����t7��t2���t-�D$P�L$Q���D$    蒣���������_^]3�[��� _��^][��� �̃�V��~(t#h(h hk2  h����  ��2�^��ËF(����   �N$���D�����   �x�   u{Sj���r���؄�tQ�T$R�D$P���D$    �����؄�t2�|$�th�h h�2  h���<�  ��j ���q����u2�h  ���n�����u2ۊ�[^���h`h hp2  h�����  ��2�^���������������̃��D$SU3�;�VW��l$�l$�l$t�(�~�L$Q�ǍT$��R�ΉF賗���؄ۉ~��   �|$�  u{�D$P�L$Q�������؄�td�T$;�|\�|$;�vR3Ƀ~2��3�;Ѝ�   r<w;�r6�T$R�Ήl$�l$�Sv���؄�t�D$ ;�t�L$�U���p����u2�_^]��[��� �����j�ha�d�    P��SUVW�  3�P�D$ d�    �ًS���T$��   ����3�C�9h�p�d:t�F;�tUP���p:�T$�n�n�n�C3�ǉ�H�H�H�H�H�H�H�KωL$�L$�l$(t	��R���T$���� ;��D$(�����T$�{����k�L$ d�    Y_^][����C    �L$ d�    Y_^][������������V��L$�F�VPR��F �    �     �@    �F �_����F����t�F^� ��������������j�h��d�    P��H  訴 �  3ĉ�$�H  SUVW�  3�P��$�H  d�    ��$I  3�;����t$�D$ �\  ���� ����  �_9�$I  u��$I  ;Gu���',�����}  ��$I  3Ƀ�2���l$��   �t��   w	��$�@  �V�j������D$����  U3�SV���}6��;��  ;���   ��$I  ��$I  PQSUV�L$T葅���3҃�2��3��|$D2Ǆ$I     ����   ��   ;��Ä�t
W�L$D�P6���L$@Q�L$$�R�����Ƅ$I  t��$I  R�L$D�%6���\$$��t=�|$( � @u3��$I  ;D$0u&��$I  ;L$4u�L$��R$�D$@P�҅��D$��D$ ��Ƅ$I  t�L$ j �Tm���L$@Ǆ$I  ����谅���D$����   P�n����D$���   W�L$$�����D$$����$I  tw�|$( � @um��$I  ;L$0u`��$I  ;T$4uS���� ��t�_ ���:�����@ �:���@ �G0 ��P$W���҅��L$ �D$Ǆ$I  ����蘚���D$���Ǆ$I  ����t
�L$ U�yl��2���$�H  d�    Y_^][��$�H  3��Ф ���H  � ������������̃�U�l$Wh�   j V���D$     �@� ����uL�D$P�L$Q��������t/�|$�� t-h�h�h�  h���`�  ��j ����k��_2�]���SV���V���؄�t3�VR���V���؄�t"�F8Pj����S���؄�t�N@Qj���lT���؃�uc�l$��|M��t�V R���]V���؃�|7��t3�F<P���b���؄�t"�N0Qj���S���؄�t�V4Rj���S����j ���&k����t��u%hhh�h�  h����  ��[_2�]��Ã~0 t�~4 u1�G��2}�F0��F<�F0   ���n���~4|�F4d���F<��[_]������j�hێd�    P���   �  3ĉ�$�   SUVW�  3�P��$  d�    ��$   ��l$�D$H�D$�L$83�Q�T$4R�͉l$0�\$8�\$@�\$D�\$H�H������D$,t�D$@����$  ��  �D$0=����  =� uG�T$<3Ƀ}2��3�;Ѝ�   ��   L|�D$8;�sBh�hth�  h���B�  ���L$(SǄ$  �����i���D$���?�����  �L$Q���D$ �P���L$���  �yN���F�������D$��  �W���w���$�   ��]��h�   �D$PSP�_� VW�t$`��������؃�����  �L$ Q3��T$ R�͉t$(�t$,�t$$薏���؄ۈ\$�8  �|$ � @�  9t$$�a  �\$ 	���R  �L$L�T$P���ĉ�L$d�P�T$h�H�P�*����;�uz�D$lP�+}������ud�L$l�U �R ���ĉ��$�   �H��$�   �H��$�   �H���҃�u,�L$L�T$P���ĉ�L$d�P�T$h�H�P�G*����;�u�0h���)����V�� �����uLh8hth;  h���z�  ����t��Pj����h�hthK  h���O�  ����  �uV�N|��������   �D$lP�9|��������   �L$�A��ti��t;����   �y���}x��/��/��/�L$l��/�T$p�D$t�L$x�O��/��/��/�T$l��/�D$p�L$t�T$x�&��/��/��/�D$l��/�L$p�T$t�D$x�L$l��T$p�V�D$t�F�L$x�N�T$\�U�D$`�E�L$d�M�T$h�U��$�   �E(�}0�    ��$�   ����� ��tRU� ����tE���   �L$L���   �T$P���   �L$T���   �T$X���   �L$|���   ��$�   ���   �t$H�T$$U���   ��$�   ��$�   PQ�L$$RS�������ǅ�       tU���d5����u�E �Pj���ҋL$(j Ǆ$  ������e���l$�;���h�hth
  h���L�  �D$' �\$'��V�L$,Ǆ$  �����e���Ë�$  d�    Y_^][��$�   3��� ��  � hlhth  �2���h(hth�  h���ѽ  ���L$(SǄ$  �����9e���D$�hhhth�  h��蚽  ��j �Q����D$SV��W�L$Q���D$j�΋ډD$�F0 �(]����t �T$SWR���&i����t�D$SWP���$���_^[� �������������̋D$S2ۅ�V��u#h�h�h�  h���	�  ��^��[� y#hXh�h�  h����  ��^��[� W�|$��$hh�h�  h��踼  ��_^��[� U�l$��}%h�h�h�  h��苼  ��]_^��[� j P�������t9�D$Pj�Ή|$�!\���؄�t�L$Qj�Ήl$�	\���؄�u���|�����]_^[� ��̃�V��2���x@  �  �F(SUW3�;�~:�N$���D�;�t,�P������t�P;׋H|;�s3�3ҋ�h���3�3��P���҉D$�|$�D$;|$w�|$ ��   ��P���D$ �|$�ҋ����t3�;�wrr;�wl3�9L$,j ���T$R�L$���y�����tM�D$;D$,t]��t?�D$ P�L$Q���֓����t*j ���b����t�|$��o����|$  u�|$$ �]�����D$�RP����_]2�[^��� _][�^��� ��j�h�d�    PQSUVW�  3�P�D$d�    ��~�5  �L$��6���|$(3�ωl$ ��c�  ����   Uh  ��������؄���  W�L$�
7���D$P���_���؄�t%�OQ����]���؄�t�T$(Rj�Ήl$0�Z���؍GP�L$��6����tR�L$Q����^���؄�t@�W,R���]���؄�t/�D$(Pj�Ήl$0�Y���؄�t�OP�T$(R�L$,j���Y���؋��������  ���  �oT���o�  ����   j h  �������؄���   �GX�L$(Qj�ΉD$0�JY���؄�th�W`�D$(Pj�ΉT$0�/Y���؄�tM�Od�T$(R�L$,j���Y���؄�t2�Gh�L$(Qj�ΉD$0��X���؄�t�Wl�D$(Pj�ΉT$0��X����U�L$�5����t�L$Q���]���؋��9�����t@��t>�Wp�B��pj ���Ѕ�t+j h  ���@����؄�t��B V���Ћ��������u2ۍL$�D$ �����r8���ËL$d�    Y_^][��� j h  �������tڋL$(V� �  ������褄����u����������������QV��~u�L$V�<������D$�D$^Y� U3�Uh  �������D$�  SW�|$V�������؋Έ\$�7�����u_[]�D$^Y� ����   �~��   ���  �Ƅ@  9n|�n�GP���Ɓ��;�~+�ߋL$���  �W�s������uW���/�����L��u�h�/������h�/������h�/������h 0�������h�/������h�/���ߑ��h�/���ӑ���F��t&�v��~� g��t��~h gjVP�� ��_[�D$]^Y� ���������̋T$VWR���"������u#h�h�hw  h���ö  ��_2�^� �~ t#h@h�h{  h��蚶  ��_2�^� �~( t#h h�h  h���q�  ��_2�^� j R���������t�~_^� ̋T$VR�������u"h�h�h�  h���&�  ��2�^� 9Ft"hph�h�  h�����  ��2�^� �~(t"h4h�h�  h���׵  ��2�^� �F(��~V�N$���D���tH9PuCSj j��������؄�t���ہ����u2ۋ��΁����u2ۋ�B���Њ�[�F    ^� h�h�h�  h���X�  ��2�^� ���������������h  �F���������h  �����������V��~th  ����^Ã~( t h�hXhd  h����  ��2�^Ã~ thhXhh  h���ƴ  ���F   �^���������V��~u-�~th 	h�h�  h��舴  ���F    �^�h  � ���^���������������h  �f���������h  �����������h  �F���������h  �����������h   �&���������h   ����������h"  ����������h"  ����������h#  �����������h#  �v���������h!  �����������h!  �V���������h%  ����������h%  �6���������h&  ����������h&  ����������h  �f���������h  �����������j�hY�d�    P���   �  3ĉ�$�   SUVW�  3�P��$�   d�    ��$�   ��L$D�D$ �A��3ۉ�$�   ��    �L$$Q�T$R�Ή\$$�\$ �\$�S�������  �D$=	  wR=  �  -  t8��t����  Sh �D$$P�L$PQ�   Sh �T$$R�D$PP�   Sh �v-  ��  -�� ��   ���j  �D$$P�L$Q�Ή\$�:������M  �|$  �?  �T$$R�D$P��蓊�����&  S���sY�����  Sj��L$$Q�T$PRS����������   �D$������   �F(;�~�N$���l��3�3���t �}  u9}u9}u��B���Ћ��3�L$,�����L$,Qj����A����tj j��T$$R�D$PPj ���b�����u���D$����tk��tg�F(��~�N$���D��3�;�uN�}  uE�} u?�} u9��B����3�;�r*w;�v$+�ϋ��׃���������wr�����w�}�M3ۋ~�σ��NS���BX�����~tv9\$t�|$ ;�ur9\$������   �L$$Q�T$R�Ή\$�~����t��|$�� u��D$$P�L$Q���������t�S����W����t�Sh�� �T$$R�D$PP�g����D$�����7h�   �T�����D$ ;�Ƅ$�   t�T$DR���"����3���D$   �L$DǄ$�   �����p?���D$��$�   d�    Y_^][��$�   3��ŏ ���   � ��h  �����������h  �V���������h  ����������h  �6���������V��~ Wth�	h�	h61  h���]�  ���|$Wh`/�kj������u#hP	h�	h91  h���+�  ��_2�^� �|$ Ut&�l$��~�|$���|��2|�~2}]_2�^� �F�n�D$Sh  ��������؄��  j h��  ���4����؄���   W����Q���؄���   j h��  ���
����؄���   �L$Qj���D$   �:N���؄�t�T$Rj���D$$    �N���؄�u���z����tO�D$P����y���؄�t0�L$Qj�Ήl$ ��M���؄�t�T$ �D$ Pj�ΉT$(��M���؋��Dz����u2ۋ��7z����u2����tj h�   ���M����؄�uh  ���{�����[]_^� ��SV��F(��~"�N$���D���t�x�   u����y�����hH
h 
h�1  h���z�  ��2�h  ��������u^[�^��[��������������V���P�҃~( t h�
h�
h�2  h���'�  ��2�^Ë�PSUW����3�Uh�  �΋��s����؄�tE�F3Ƀ�2��3҃�2��   ��   �D3���QP���WZ���Ί���x����u2ۋ�B����_]��[^���������SU�l$W���������D$Pj���b<���؄�tC�L$VQ�������3�9t$~%��$    ��tW����?������2����;t$��|�^_]��[� _]��[� ̋D$��V��t
P�  ^� j h� ������tCSj h�� ���l����؄�th`/���*O���Ί��!x����u2ۋ��x����u[^� ��[^� ���̃�\�  3ĉD$XVW�|$h��~�|$}_�^�L$X3�苋 ��\� SU�o����  ����$    ��|$����  �E �P8���҅���  ��|@   uV���q#�������m  �Eh`/P�(g�������T  ;��   �H  �E ����ҋ����5  ��Hg�)  �����  �D$P���*� ��L$X�P�T$\�H�L$`�P�D$Xh`/P�T$l�f��������  �L$(Q�Hg�F��P�T$\R�f��������  �D$8P����!��P�L$\Q�ff��������  �T$HR�������P�D$\P�Af�������m  �~uh g�MQ���@  �,�����K  �EP�f������t$�����Ph�h�  h���8�  ���  U�j� ���͋��n� ��u)����   h�hXh�  h��詩  ����  ��u!hhXh�  h��脩  ���  ��|@   ��  ���   ����  ��~	��2��  ���   Rt��y  ��2|
�~2�j  j h� �������؄��R  jj��� P��j h�� ���r����؄��"  �T$XR���,L���؄���   �EP���L���؄���   �E(�L$Qj�ΉD$�xH���؄�t{�U0Rj���J���؄�th�EP����K���؄�tW������P�t����t���   ��F�L$Qj�ΉD$� H������t���   ��F��t�T$Rj�ΉD$��G���؋��pt����tT��tRj h � @�������؄�t>��t�~ ���f�����@ �[���@ �F0 �E �P V���҅������t����u2ۋ��t����u2ۋ��   ���K����L$h]��[_^3�複 ��\� ���̃�@�  3ĉD$<�D$DS�U�D$ 3�3��y2V��W�T$R�L$�l$�l$ ��   �����D$P�l$4�l$8�l$(�l$,3�������u3�_^][�L$<3��%� ��@� �|$� t!h�h�hh  h����  ���  �L$���;�+|�T$;�s!hXh�hm  h���ʦ  ���r  �|$�D$,P�L$Q���=����;��T  �|$�� thh�h{  h����  ���;�|$,u9l$0th�h�h�  h���T�  ����T$<R���8����u3�U���M������  ;���  �D$<h`/P�6a������u�p�  ;�tN�����ЍL$,��Q�����P�T$@R�b������uPhhh�h�  h���¥  ���   �g  �L$<�T$@���ĉ�L$T�P�T$X�H�P� ������;�u&h h�h�  h���>�  ���   �  �D$ P�L$Q�L$��}����;���   �|$�� t#h�h�h�  h��� �  ��3��   9l$$(|9l$ w hxh�h�  h����  ��3��t;�u-��������;�u h8h�h�  h��辤  ��3��C��D$�R$P���ҋ�;�u)h h�h�  h��芤  ��P��j������D$(��L$U��K����t;�t;�t�L$S�$�����u3��L$U��K����u3��L$L_��^][3��'� ��@� ������̃�<�  3ĉD$8SUV��2���x@  W�  ��P�ҋЋF(3�;ŉT$�6  �N$���L�;��$  �A���Шu3h�h�h�  h��謣  ��_^]2�[�L$83�蒃 ��<� 9i:|9is3hph�h�  h���m�  ��_^]2�[�L$83��S� ��<� �y;�rjw;�rd�����;�wWr9D$wO�L$+ˋ��RQ������؄�t�L$PQ��������؄�u�T$UR�����_^]��[�L$83���� ��<� hh�h�  h���Ǣ  �L$X��_^][3�2�譂 ��<� �F�3�;��#��BW���Њ؄�u;�v��BU��3��Њ�3��ۉD$$�D$(�D$,�D$0�D$4�D$8�D$<�D$@�D$D�N����L$$Qj ����(���؄��6���j�T$(h��R�U� �����Ä�uC;�v7��PU��3��҄�t�D$$Pj ���(��j�L$(h��Q�� �����Ä������;~t�~����T$�D$�D$R�D$P�Ήl$��o���؄�������|$u9l$�}���|
9l$�q���2��������̃�UVW�|$ W��������u'h�hxh�  h���O�  ��_^2�]��� �~ t'h0hxh�  h���"�  ��_^2�]��� �~( t'h�hxh�  h�����  ��_^2�]��� �F��S'��  t,��Pj ���҄��Ê�[_�n^]��� ��  u��[_^2�]��� 3������L$�D$�D$�D$PQ���n���؄�t<�D$;��b  ��  u2ۊ�[_^]��� ��  u�~�����   ��n��[_^]��� ��  u	�~|l��؁�   u	�~�l��ǁ�!  u	�~6��북�"  u	�~&��륁�#  u	�~�o�딁�%  u	�~���냁�&  u�~\���o���="  �D$$uz��!  ur�~ul�~���|c�T$R�D$P���D$    �
x����tF�|$"  u�D$$ j ����F����t*�|$$ u#�L$Q�T$R���D$    �Jm���|$!  t&h�hxh=  h����  ��W��������؄�������D$�L$Q�T$R�ΉD$�yw���؄������9|$�����hHhxhG  h��輞  ��j ��2��.F����[_^]��� ��Vh  ��������uQ�`/�d/j j(���ĉ�h/h��  h  �P�l/�Hj j �ΉP������th  ������^������������̃�V��h  �F    ������uX�D$P��9����j j���̉�P�Q�P�@hP�  h  �Qj �Aj ���R����t%h  ���B���^��Ã~uh @ �������^������̃�V��   9Ftah  ������uS�D$P��z�#���j j���̉�P�Q�P�@hs�  h  �Qj �Aj �������th  ������^������������̃�V��~�^���h  ������uS�D$P�0�����j j���̉�P�Q�P�@ht�  h  �Qj �Aj ���<����th  ���,���^���������̃�V��~�^���h   ������uS�D$P��� ���j j���̉�P�Q�P�@hu�  h   �Qj �Aj �������th   ������^���������̃�V��~�^���h"  ������u\�~"��|S�D$P� y�
���j j���̉�P�Q�P�@hw�  h"  �Qj �Aj ���3����th"  ���#���^����������������̃�V��~|o�~�o�|fh#  �������uZ�D$P�0v�
���j j���̉�P�Q�P�@hx�  h#  �Qj �Aj �������th#  ������^��ð^����������������̃�V��~�^���h!  �c�����uS�D$P��F�	���j j���̉�P�Q�P�@hv�  h!  �Qj �Aj �������th!  ������^���������̃�V��~|r�~���|ih%  �������u]�D$P�PU�����j h�  ���̉�P�Q�P�@hz�  h%  �Qj �Aj �������th%  ������^��ð^�������������̃�V��~|o�~\��|fh&  �Q�����uZ�D$P� w�n���j jt���̉�P�Q�P�@h{�  h&  �Qj �Aj ���
����th&  �������^��ð^����������������̃�V��h  �F    �������uS�D$P��S�����j jr���̉�P�Q�P�@h@�  h  �Qj �Aj �������th  ���r���^���������������̃�Vh  ���P�����uS�D$P��R�m���j j���̉�P�Q�P�@h`�  h  �Qj �Aj ���	����th  �������^�������V��h  �F    �������uQ�`/�d/j j���ĉ�h/hp�  h  �P�l/�Hj j �ΉP�����th  ������^������S�\$WS���T������t_2�[� �L$��~��D$= ��|�V�t$�>�   u�~ t�~ tPQjS���+�����u^_2�[� �F�NPQ���0���ϊ��������u2�^_��[� ��������̃��D$��UVW���D$ t�  �l$,��t�E     �|$0��t�    �~u_^2�]��� Sh  �����؄���  �D$P�L$Q���D$    �o���؄���  ���  9|$t!hPh(h�1  h���Ζ  ���  �T$(R���*)���؋F(��~�N$���L��3Ʉ��y  �~n���l  ���d  9y�[  �����3Ƀ~2������   ��-��3�;��5  w;��+  3��T$2ۅ҉|$�|$u!h��hX�h�  h��� �  ���k  �D$��u!h��hX�h�  h�����  ���B  �L$Q�T$,R�Ή|$�|$ �|$0�|$$�|$(��c�����  9l$(t#hP�hX�h�  h��覕  ��2���   9|$ ,|�|$s#h�hX�h�  h���t�  ��2��   �D$P�L$,Q�Ή|$0�|$$�|$(��m���؄���   9l$(uf9|$ |`�|$rW�T$Rj��� %���؄�ta�|$}h��hX�h�  �:�D$Pj����$���؄�t59|$}7h��hX�h�  �h0�hX�h�  h��辔  ��2�W���1<���l$0����   �L$03�Q���D$�D$4�|$,�|$ �53���؄�tO�D$,;�t�T$0��D$(Pj���C$���؄�t-;�t�L$(�M �T$Rj���$$���؄�t�D$4;�t�L$�W���;����u2�j ���;�����|$4u2ۄ��D$    tH�T$R�D$P���l���؄�t1�|$�   t7h�h(h#2  h���ɓ  ��j ���=;��2�h  ����c����t@�|$ u9�F��2}��t�E ��t&�N��[�_^]��� ��t�E    ��t�d����[_^]��� ���������������SU�l$VW�|$����|��u3��D$Pj�|$��2��3���~����t�L� Q���������;�|�_^][� ��j�hݏd�    P���  �  3ĉ�$�  SUVW�  3�P��$�  d�    ��$  �������҅�u#h�h�h�  h��藒  ��2��  ��$  Q���.�����$�  �H��$�  �P��$�  �@�   9o��$�  ��   V�3!�������2  V���������!  �L$���������   j ���D$ �$P��Ǆ$      �҅�t'�D$P��������L$��Ǆ$   �����B����  �L$Ǆ$   �����)�����  ��B(����=   @��  V�E����؃�����  ���A?����u���D��;�|��BXj ���Ћ��u+j ���X������u��PP���$P���pP ����]  �U �B(����=   @�<  U��������U �؋Bj�����!  V�P< ����t~V��  ����uq�L$能  �����   ���D$�$P��Ǆ$     �҅�t'�D$P�������L$��Ǆ$   ������  �  �L$Ǆ$   ������  �����V�E! ������������� �����������$�H
�L$T�׍ �L$TQ�Ή�$  �D; �T$TR���(����L$T��Ǆ$   ����� �(  �L$T�� �D$TP��Ǆ$     �-C �L$TQ��������L$T��Ǆ$   �����ۍ ��  �L$T�}� �T$TR��Ǆ$     �: �D$TP�������L$T��Ǆ$   �����d� �  �L$T�֏ �L$TQ��Ǆ$     �o: �T$TR���S����L$T��Ǆ$   ����轏 �S  ��$$  �܍ ��$$  P��Ǆ$     ��E ��$$  Q��������$$  ��Ǆ$   �����
� �   �U �Bj����j h� ���;����؄���   j h�� ���#����؄���   ��$�  Q����1���ϊ���Z����u2��x��ttj h�� ��������؄�t`��B W���Ѕ��Ä�uh�h�hD  h���E�  �����{Z����u2��"��t��|@   u�������t
V���S�����j h�����s�����t���8Z����u2ۋ��+Z����u2ۊË�$�  d�    Y_^][��$�  3��m ���  � ��
�
�
:
:
�
�
�����������̋D$��u!hDh$h(  h���o�  ��3�� �     �D$�����������̋D$�T$R�D$����� �����������V��2��~tt�F(��~H�N$���D���t:�x  u1j h��  ���i�����tD�T$SR��������Ί��Y����u'[^� h�h�h
  h��轌  ��2�^� ��[^� ������������̃�SUVW�|$ 3�;���t�/3��{��   �D$P�L$Q�ˉl$��d������   �D$=��  uz�T$R�ˉt$������t1�|$W�Iq ������u��t��Pj������   ���|$ uh h hI  h�����  ����t�7�2��t.��Pj�����!���th h hR  h��迋  ��j ���33��_^��][��� �������j�h�d�    PQSVW�  3�P�D$d�    ��2ۃ~th(hhu  h���Y�  ���~�[  �~( t3h�hh{  h���-�  ��2��L$d�    Y_^[��� �|$$����K��P�L$(����L$$�D$    �]������   j h @ ���G����؄���   j h @ ���/����؄�t�D$$P���]/���؋���V����to��tm�L$Q���K�������Ph @���������Ί��V����t>��t<���tK����t�   ����RK�������Ph3 @��������Ί��uV����u2�j j���������u2ۋ��WV����u2ۋ��JV����u2ۍL$$�D$������	���k�F(��~F�V$���D���t8�x  u/j hP�  ���5����؄�t9�D$$P�������Ί���U����u �h`hh�  h��苉  ��2ۊËL$d�    Y_^[��� ��������������̃�U�l$��V��u
^3�]��� �E     �~th�h�h�  h���!�  ��W3��~�|$u�D$P���t���|$�   �L$Q�T$R�Ή|$ �wa������   �D$=P�  SuG�D$P�Ή|$ �3�����t"�\$S��G��������uA��t��Bj����hlh�h�  ����thlh�h�  h���n�  ��j ����/��[��th`/���m��3��} ��_^��]��� ��������������V��~
th�hlh�  h����  ���F(��~H�N$���D���t:�x  u1j hs�  ���O�����tD�T$SR��������Ί��T����u'[^� hhlh�  h��裇  ��2�^� ��[^� ��̃�U�l$��V��u
^3�]��� �E     �~t�~
th0hh   h���K�  ���~���|�S�D$P�L$Q���D$     3��_����t~�D$=s�  WuG�T$R�Ή\$ �s�����t"�|$W��� �؃���uA��t��Pj����h�hh4  ����th�hh8  h��讆  ��j ���".��_3��] ��[^��]��� ��������������V��~th�h�h\  h���^�  ���F(��~H�N$���D���t:�x  u1j ht�  ��������tD�T$SR�������Ί��UR����u'[^� h�h�hi  h����  ��2�^� ��[^� ��̃�U�l$��V��u
^3�]��� �E     �~~�~th�hph�  h��蛅  ���~|l�|�W�D$P�L$Q���D$     3��^����t~�D$=t�  SuG�T$R�Ή|$ �������t"�\$S�L ������uA��t��Pj����h8hph�  ����th8hph�  h�����  ��j ���r,��[3��} ��_^��]��� ��������������V��~th`h<h�  h��讄  ���F(��~H�N$���D���t:�x   u1j hu�  ���������tD�T$SR���n����Ί��P����u'[^� h�h<h�  h���C�  ��2�^� ��[^� ��̃�U�l$��V��u
^3�]��� �E     �~~�~thh�h   h����  ���~�l�|�W�D$P�L$Q3��Ή|$ �W\����t~�D$=u�  SuG�T$R�Ή|$ ������t"�\$S�X ������uA��t��Pj����h�h�h1   ����th�h�h5   h���R�  ��j ����*��[3��} ��_^��]��� ��V��~th�h�hY   h����  ���F(��~H�N$���D���t:�x"  u1j hw�  ���O�����tD�T$SR��������Ί��O����u'[^� hhh�hz   h��裂  ��2�^� ��[^� ���j�hK�d�    P��SVW�  3�P�D$d�    ���\$,��u3��L$d�    Y_^[��� �    �~݃th�h�h�   h����  ���&��|��D$P�L$Q���D$    3��Z������   �D$=w�  ��   �"��}[j8�0&�����D$���t$$t���z� ���3���B$W���D$(�����Ѕ���   ��Bj����hHh�3�h�   �[�L$Q�ωt$�������t"�\$S�޸ ������uA��t��Bj����hlh�h�   ����thHh�h�   h����  ��j ���(���\$,3����3���L$d�    Y_^[��� ���������V��~th�hth!  h��辀  ���F(��~H�N$���D���t:�x#  u1j hx�  ���������tD�T$SR���~����Ί��L����u'[^� hhth!  h���S�  ��2�^� ��[^� ��̋D$��SV3�;Ƌ��  �0�{��   �{�o���   �{thHh hS!  h����  ��U�D$P�L$Q�ˉt$����gX������   �D$=x�  uZ�T$R�ˉt$�$�����t5W�|$W�El ������u��t��Pj������D$ �0�   ��_u6h�h hm!  ����u3��h�h hw!  h���H  ��j ���&����u�����]^[��� ^3�[��� V��~th@hh�!  h����~  ���F(��~H�N$���D���t:�x!  u1j hv�  ���?�����tD�T$SR�������Ί���J����u'[^� h�hh�!  h���~  ��2�^� ��[^� ��̃�U�l$��V��u
^3�]��� �E     �~~�~th h�h�!  h���;~  ���~6��|�W�D$P�L$Q���D$     3��V����t~�D$=v�  SuG�T$R�Ή|$ �c�����t"�\$S�����������uA��t��Pj����h�h�h�!  ����th�h�h�!  h���}  ��j ���%��[3��} ��_^��]��� ��������������SV��2ۃ~th h�h!"  h���K}  ���F(��~G�N$���D���t9�x%  u0j hz�  ��茿����t<�T$R�������Ί��CI����u!^[� h�h�h'"  h����|  ����^[� ������̃�SU�l$V3�;����   �u �{�t$��   �{�����   �D$P�L$Q���D$$�����U������   �D$=z�  uZ�T$R�ˉt$�������t5W�|$W�����������u��t��Pj������u �D$    ��_u8h� hh h�"  ����u�t$�h� hh h�"  h����{  ��j ���f#����u�D$�����D$^][��� ^]3�[��� ��SV��2ۃ~thh!h@!h�"  h���{  ���F(��~G�N$���D���t9�x&  u0j h{�  ���ܽ����t<�T$R���\����Ί��G����u!^[� h� h@!h�"  h���1{  ����^[� ������̃�S�\$W���    ��D$    ��   �\����   U�D$P�L$Q�σ���kS������   �D$={�  uY�T$R���D$    �$�����t+V�t$V��z �����u��t��Pj������   ^�; u6h�!h�!h#  ����u3��h�!h�!h#  h���Mz  ��j ����!����u�����]_[��� _3�[��� �����SV��2ۃ~th�"h�"hB#  h����y  ���F(��~G�N$���D���t9�x  u0j h@�  ���<�����t<�T$R�������Ί���E����u!^[� h0"h�"hH#  h���y  ����^[� ������̃�UVW�|$3�;���u_^3�]��� �7�}�t$uW����_^�D$]��� �D$P�L$Q���D$$�����Q������   �D$=@�  uY�T$R�͉t$�x�����t4S�\$S����������u��t��Pj�����
�7�D$    ��[u8h#h�"h�%  ����u�t$�h#h�"h�%  h���x  ��j ��� ����u�D$�����D$_^]��� ������SW��2ۃth�#h�#h�%  h���Kx  ���G(���3  �O$���D����!  �x  �  j h`�  ��耺�����  �T$R��������؄���   V�t$����   j ha� ���G����؄���   ��P W���҅�������C����tw��tu��|@   u���?�����ta�|[����  ��tPj hb  �������؄�t<V�������؄�t!j h�����ʹ���؄�t���C����u2ۋ��C����u2�^j ho  ���蛹����t���`C����u2ۋ��SC����u!_[� h`#h�#h&  h����v  ����_[� ������̃�SUVW�|$ ����t���xs���t$�����u_^]3�[��� �    �{t(hx$hT$h�&  h���v  ��_^��][��� �{uWV����n��_^��][��� �D$P�L$ Q���D$$    ��N�����'  �D$=`�  ��   �T$R���D$     ������t �|$W谼������u0��t��Pj����h$hT$h�&  h����u  ���   ��   ���D$P�L$ Q���D$$    �GN������   �t$��a� u;�L$ ��tU��B$S�Ѕ��D���th$hT$h�&  h���qu  ���I3��E��b  u�|$  t�L$ Q��������u���j �������t��o  �t���X�������j �����_^��][��� ��������������j�hx�d�    P��$SUVW�  3�P�D$8d�    ��2ۃ	th8%h%h�&  h���t  ���G���t$H��   ��P(���҃���   V�{U �����D$Htx���y���3����D$���  3퍤$    ����  �D$H�@�P�L$�����L$LQ�T$R���D$H    �,����L$���D$@������������;t$|��  �G(����  �O$���D����q  �x  �d  ��B����j hp�  ���7����؄��'  ��B(����Phq  ���������t����?��V�������؄���   �t$L����   j hr� �������؄���   ��B W���Ѕ������?����tw��tu��|@   u���������ta�|[����  ��tPj hs  ��腵���؄�t<V���G����؄�t!j h�����c����؄�t���&?����u2ۋ��?����u2�j h  ����5�����t����>����u2ۋ���>����u2ۋ�B���Є�u 2��h�$h%hG'  h���}r  ���ËL$8d�    Y_^][��0� �̃�SUVW�|$0�������t����n���t$,��u_^]3�[��� �D$4���    u����{uPWV���Ф��_^��][��� �D$P�L$4Q���D$8    �{J������   �D$0=p�  ��   �T$R�D$4P���SJ������   �|$0q  �th�%h�%h�0  h���q  ��j �����V���������t
��uu�h�s�   �L$Q�T$4R���D$8    ��I����tN�D$0=r� uf����   ��P$S���҅���   ����   ���t;h|%h�%h�0  h���q  �����j ���y����u���_^��][��� 3���=s  ud��t`W��蟭����u����O�D$P��W�g���P�������P����������t)���    ���   �����   R���ғ����Pj����j ��������u����|$0  ��W�����������I�������������̃�SUV�t$�FW3�;ǋ�t�N��QWP�T ���T$Rj�͉~������؄�t�D$P���E���9|$�|$_^]��[��� 3��L$Q�͉|$�-����|$���Ä�t:W��.�������D$t)�T$R���"���D$��;D$�D$|�_^]��[��� ��t��Pj����_^]2�[��� �����������+� �����������QV�t$��u�D$���^Y�W�|$����   �dX���%  �=hX ��   �f���΋�v+����I f=� s�f��vf=� s�A����f��w�f�9 ��   f�: ��   V�L$����W�L$����j��L$�z���Pj��L$�n���P�dXh  P�@!���L$u�N����L$�E���_���^YÃ�u�4����L$�+���_3�^YÃ�u�����L$����_�   ^Y������L$�����WV�� ��_^Y�j�Wj�Vh  P�D!��t���t���t�WV跋 ��_^Y����������������ߌ �����������鼍 ����������̸��������������[����������������������������̋D$����   �$� ?
�   ø   ø   ø   ø   ø   ø   ø   ø   ø   ø   ø   ø   ø   ø   ø	   ø   ø
   ø   ø   ø   ø   ø   ø   ø   �3�ÍI ?
�>
�>
�>
�>
�>
�>
�>
�>
�>
�>
?
�>
�>
�>
�>
�>
�>
�>
�>
�>
�>
�>
?
?
?
�������̃�t&��t!��t��	t��t��
t��t��t3�ø   ������������������D$�L$��;���  ����  �Q�����  �������  �$��D
Q��j������� {���Q��j�������@<���Q��j��������'��Ë��؃�����   ���  ���  ��������Qtj�N����5H'���j�=�����'��Ë��؃�����   ����   ���������Qtj�����5@'���j������p&����؋���������Qtj������58'���j�������'��ÍA�����   �$��D
�����K������0'�������'�������'�������'�������'����������'������p&�������'�������'������@<������('������ '������'������'Ë�����������  Q��j������5'���Q��j���������'���Q��j��������'����؋����d�����Qtj�����5 '���j������'���Q��j���q�����'���Q��j���[����0'���Q��j���E�����'���Q��j���/�����'��ÍA��؃���   �$�`E
����&�����&�����&����H'����@'����8'����'�����&�����&���� '�����&�����&�����������+�����&�����&�����&�Q��j�m����'��Ã�
����t��tQj�M����h�����pD���&Ë��؃�	��t��tQj�����P'�����&����Ã�	����u��&Ë�������Qtj������h�����&�j�������&���Q��j�������5�����Q��j�������5�+���Q��j��������&���Q��j���s�����&���Q��j���]����x&���Q��j���G����p&�����Ë�8@
N@
�@
A
!B
B
�B
�B
mC
�C
�D
@
"@
�@
�A
B
SB
iB
�C
D
%D
;D
QD
gD
}D
>A
IA
TA
jA
�A
�A
�A
�A
�A
�A
�A
(A
3A
_A
mA
xA
�A
�A
�A
�A
�A
�A
�A
�A
�A
�B
�B
�B
�B
C
@A
KA
�D
>C
PC
YC
�B
�B
�B
�B
C
C
#C
GC
,C
5C
�����������̋L$3�+�t��t��u�   ø   �3��������������̋L$3���w3�$�0F
3�ø   ø   ø   ø   ø   ø   ø   ÐF
F
F
F
F
F
F
F
F
F
F
#F
)F
�����������̋L$3���w-�$��F
3�ø   ø   ø   ø	   ø   ø   ÍI �F
�F
�F
�F
�F
�F
�F
�F
�F
�F
�F
�F
�F
�L$3���t	��u	�Aø   ������̋L$3���w�$�(G
3�ø   ø   ø   ÐG
G
G
!G
�������̋D$�� t��t��u�   ø   �3���������������̋L$3�+�t��t��u�   ø   �3��������������̋L$3���w?�$��G
3�ø   ø   ø   ø   ø   ø	   ø
   ø   ø   Ð�G
�G
�G
�G
�G
�G
�G
�G
�G
�G
�G
�G
�G
�L$���3���w�$�PH
�   ø   ø   ø   ÍI 5H
;H
AH
GH
�D$�� t��t��u�   ø   �3���������������̋D$��w ���H
�$��H
�   ø   ø   �3�ùH
�H
�H
�H
�H
 ������̋L$3���w9�$�8I
3�ø   ø   ø   ø   ø   ø   ø   ø   ÍI I
I
I
I
I
I
#I
)I
/I
���̋��     �@    �SU��V�u 3�;�t���F;�t	P�6r ���6;�u�u;�] t&W���G;Ë6tP�!�����_W�!����;�u�_^�]][����S�\$U3��W��v5Vj� ��������tS� ���F�O����w^_][� ^_��][� _��][� ����SUW�|$��3����v5Vj�E ��������tW�6 ���F�K����s^_][� ^_��][� _��][� SUW�|$���3����v5Vj����������tW�����F�K����s^_][� ^_��][� _��][� �������������̋D$SU�ًL$PQ�m��������t8VWj3����������tj�y�����w�S����{���n_�3��^][� ��������;��������������j�h�d�    PQV�  3�P�D$d�    ��t$�T'�N0�D$   �R����N,�D$�E����N(�D$�8����N$�D$�+����N �D$�����N�D$�����N�D$�����N�D$������N�D$ ������N�D$����������L$d�    Y^������������j�hP�d�    P��SUVW�  3�P�D$ d�    ���D$0�wP������h�f�L$Q������V�T$43�R�ȉ\$0�t����oP���D$,�T����L$0�\$(�G�������L$�\$(�7���h�f�D$P���f���V�L$4Q���D$0   �!����oP���D$,�����L$0�D$(������L$�\$(�����h�f�T$ R������V�L$Q���D$0   �����P�O�D$,�����L$�D$(�����L$�\$(�����L$ d�    Y_^][��� �j�h��d�    P��SUVW�  3�P�D$ d�    ���D$0�w P���x���h�f�L$Q���w���V�T$43�R�ȉ\$0�4����o$P���D$,�����L$0�\$(��������L$�\$(�����h�f�D$P���&���V�L$4Q���D$0   ������o(P���D$,������L$0�D$(�����L$�\$(����h�f�T$ R�������V�L$Q���D$0   ����P�O,�D$,�r����L$�D$(�d����L$�\$(�W����L$ d�    Y_^][��� �W���G8��~ V3���~S�_j ��������;w8|�[^_�h`'�O����_��������V��W�~���r����v8���   ;Ƌ�|+�P�h���_^�_^������������������́�  �  3ĉ�$  ��$  ��V��$  �D$ �  ��$  QP�T$h�  R��������|$ Ƅ$   ��   SW�|$�|$��U��I �;
ui�~4 � t3�n���h�����t%j �������8 t�>�̓��J���P����Ћ|$�? t
��BW���Ћ�Bh�&���ЍK�F4   �L$�����; u��? tF�~4 t/�n���������t!j �������8 t��̓�������P���ҋ�PW�����F4    ]_[��$  ^3��; ��  ������̋T$��t9�: t4�A��t�T$���a���A��tPR��| ��� Rh,+�| ��� ������������j�hȑd�    PVW�  3�P�D$d�    ��N��t�D$P�;���L$d�    Y_^��� �L$Q�L$ �I����>�L$�D$    �����WP���ҍL$�D$���������L$d�    Y_^��� ����������D$V�5������Dzhd'��V������^� ���N�$�z���PV������^� ������������V��h KV�b����D$�@���\$�N� �$�7���PV�@���h�)V�5����� ^� ��������������VW��h KV�����|$��W�����r����t!ht'V�������h�)V�������_^� �G���\$�N�G�\$��$����PV������ h�)V������_^� ���������������V��h�'V�����D$�@���\$�N� �$�W���PV�`���h�'V�U����� ^� ��������������VW��h�'V�1����|$��W�x���q����t!h�'V������h�'V������_^� �G���\$�N�G�\$��$�����PV������� h�'V�������_^� ���������������U�������4SV�uW�������$�������th�'W������_^[��]� ���N�����th�'W�_�����_^[��]� j ���z���j �ΉD$@�_�j����@���$j ���X����@���$j ���F����@�D$L���\$��� �$�����PW�����h�&W�������0j������j�ΉD$@�����@���$j��������@���$j��������@�L$L���\$����$����PW����h�&W������0j������j�ΉD$@�����@���$j�������@���$j���t����@�T$L���\$����$����PW�#���h�&W������0j���<���j�ΉD$@�/����@���$j�������@���$j�������@�D$L���\$��� �$����PW����h�&W������0_^[��]� ��̋D$�Pf��uKf�x�uC�x�u=�x	�u78P
u2�xu,�xru&�x�u �x8u�xxu� Ph�'Q�N������ V�pV�pV�pV�pV�pV�p
V�p	V�pV�p� V��RPh�'Q������4^� �V��L$������tf�8 t
�P�B����^� ������������V�t$W������������uh((W������_^� �������P�������P�������Ph(W������_^� ��������������U����j�h��d�    P��hSVW�  3�P�D$xd�    ��hk4�L$ �4����E��Ǆ$�       t�8 t
P�L$ �c����}��t�E���D$ ��M�L$ �} �]u�L$����Ph)���u�L$����Ph )V��������} �D$$    ��  �U�������3��(����Ƀ�4��)�L$,��    �D$(�L$0���D$(�T$$PR�L$$�-���Ph�(V�a�������N�$�A���PV�J����   ��9|$ ~,h�fV�1������N�$����PV��������;|$ |ԋD$,Ph�(V� ������} ��   �M����������D��   ��h�(��V�T$D��\$<������D$<�N�$����PV�����   ��9}~9����h�f�L$@V�\$<�����D$<�N�$�k���PV�t�������;}|�h�)V�^��������h�&V�L����D$,\$8����;E�D$$������L$Ǆ$�   ����������L$xd�    Y_^[��]� �������́�  �  3ĉ�$  S��$,  ��VW��$0  �L$t�; u�0)3�9�$   ~`U��$,  ���VS�D$h()P�YB ��$@  ��$8  ���L$Q��$$  WR��$(  PQ�L$$R��������;�$$  |�]��$  _^[3��72 ��  �  ����QS�\$��UVW���|$uh�)W�"������t$��}h�)W�������l$;�}h�)W�����������   ;���   ����   UV被 hh)3�W��t$0����������   �d$ �N;Ϳ   }�T��������Dz������;�|��u��D$W���$VhT)P�j������-��L$ �$ˋT$���$W����$Vh8)R�;����� �t$ �;��z���_^][Y� ��V���H����D$t	V�[�������^� ��j�h��d�    PQV�  3�P�D$d�    ��t$�D$hk4�N�T'�F    �F�����N�D$    ������N�D$������N�D$�����N�D$�����N �D$�����N$�D$�����N(�D$�����N,�D$�|����N0�D$�o���h�)���D$	�F4   �F8    �`���h�)�������ƋL$d�    Y^��� ��������������̸�X����������̋A(�������������VW�|$W��貿���������W�N貞��_��^� ����������V�������D$�L$PQ�N覞����^� ���������������VW�|$j ��j���]�������t2�FP����������t �NQ����������t�V(R���g�����_^� ��������������̃�VW�|$��D$P�L$Q���D$    �D$    ��������t9�|$u2�VR����������t �FP���	�������t��(V���������_^��� �����������̃��� ��������3�� �����������������$�� ��������������̃��� ��������V��N�� ��}3�^Ë�Pj ���������^���������̋D$�D$��   � �������������̃�SVW���L$�oa���w��3ۅ���   �v���3�U�I �G�,�l$�l�l$�l�l$�l�l$�l�l$ �l�l$$�,�,�l�l�l�l�l�l�l�l�l�l�G�l$(�l$�h�l$�h�l$�h�l$ �h�l$$��������;މh�^���]_^[��������̋A��~�I�D���3���������������̋A��3҅�~#V�I �q�փ��ƃ�;��\���q�\�|�^�V�t$��th�X��������t��^�3�^����������������V��������N�IN$��$��^�������̋T$V��FP�F�@���QR�BI �V �N��Q�RP�.I ��(VjP�"I ��$^� �����������VW�|$��;�t'W�.����GP�N�����V�R�N�GP�ҋG(�F(_��^� ������SV��W�~�N�0� �L$�T$��3�9D$��PQR���C_��P�F(jSj P贴 �� _^��[� ��������SVW���_����� ������   ;w ��   ������$�N� ��u$�D$��th�*P�G������?I  _^��[� �   ;�~#�W����$    �B������t@����;�|�(��|	����   �D$��tWh�*P���������H  _^��[� �T$��t+�G�ȍȃ��$Q�@����$���Qhp*R������ �H  _^��[� �D$��tB��V}h@*P�z������rH  _^��[� �O Qh�)P�Z������RH  _^��[� _^�   [� ��������������U����j�h��d�    P��hSVW�  3�P�D$xd�    ����Ph�L$4Q����j�L$8Ǆ$�       �>V��j �L$8���1V����]���\$� �$h+S�������O3��� ��~P�t$0Vh+S�����GD$<��P���b����O����$h+S�k����D$@���O���� ;�|��L$4Ǆ$�   �����p� �L$xd�    Y_^[��]� �����������j�h��d�    PQVW�  3�P�D$d�    ���D$    �|$ ���D$    �0U���N�D$    �D$   �(� �ȃ�|*�F�D�������Au�v�D�����\$����$��f���ǋL$d�    Y_^��� �U����j�h0�d�    P��hSVW�  3�P�D$xd�    ��^ ���3�����   �N��E��������D�Ez��������Dz�ٿ   ����   ������A��   ��Ph�L$4Q�����E���\$�L$4�E��$�   �$�i���E�F��N�E�   ;���Ƅ$�   ~<�d$ �V�������L$<�$�D$(�TT�����L$,�$�T���D$ ���;�|ȍL$$�   Ƅ$�    蒢 �L$4Ǆ$�   �����~� ���g����ǋL$xd�    Y_^[��]� VW�|$�G�������   9~(S��/  U�*������N��   ��~q�V��5����D{_��3���|6�Q���3����<�    �n�T(�n�T((�n�T(@�n�T(X��`��u�;�}����+ϋV�T����u���]��[_�F(   ^� _2�^� ����   �V��5��������D{i�B������Dz_��3���|6�Q���3����<�    �n�T(�n�T((�n�T(@�n�T(X��`��u�;�}����+ϋV�T����u����F(   ]��[_^� ���������V��W�N3��"� ��| �N�T$���PQR�H. ���G_^� ��_^� ������j�hX�d�    P��,SVW�  3�P�D$<d�    ��L$3�3��;����F(�D$�F���\$D�\$�D$    �D$$|>�F�D$L�N�T$�D$8+������D$0���   �L$,���L$�$�Ћ��\$8�\$,�L$�D$D�����I����ǋL$<d�    Y_^[��8� ��QSUVW�|$3�;��L$t9G|�G�t$;�t9F|�F�Y����� ���|-��t
��PS���҅�t�L$��P��Q����_^��][Y� _^]3�[Y� �������������j�h��d�    P��,SVW�  3�P�D$<d�    ��L$3�3�������N���F(�\$D�D$�\$�D$    �L$$|V�D$P�����$u�D$TP�������7�F�N�T$T�D$@+������D$8�D$�L$4R���   �L$�҉\$8�\$,���L$�D$D���������ǋL$<d�    Y_^[��8� ����������j�h��d�    P��,SVW�  3�P�D$<d�    ��L$3�3������F(�D$�F���\$D�\$�D$    �D$$|<�F�D$P�N�T$L�D$8+������$���L$4R�L$�D$<�f������\$8�\$,�L$�D$D�����+����ǋL$<d�    Y_^[��8� ����U����j�h�d�    P��(  SVW�  3�P��$8  d�    ���O�D$+ 菽 �؅ۉ\$H�,  �E�]����D�  ��Ph�L$,Q�����E�EǄ$@      ��������   ��j �L$0���uN��� �]����Auj �L$0�^N��� �]j�L$0�NN��� �E��������Auj�؍L$0�1N��� �U�E��������   �؍L$,��Ǆ$@  �����Ԝ 2���$8  d�    Y_^[��]�0 ������A��   ��j �L$0����M��� �]����Auj �L$0�M��� �]j�L$0�M��� �E��������Auj�؍L$0�M��� �U�E������u2�ٍL$,��Ǆ$@  �����1� 2���$8  d�    Y_^[��]�0 ��������D��  ��$�   �\T����$�   �PT���L$L�GT���L$|�>T���L$d�5T����$�   �)T���E$��t�     �EP�������V�u�X��������D$<��  ����  �E�E ��ݜ$�   �E�D$D   ݜ$�   t��3ۃ  ~�w�3��O�� �ESj ���$VPj�� �O���������@�����@� ������4�E�E��������   ���T��L�����z~���������zw�����������Azj�O����� �] �N;�}I�W�D�3�;��]t��D$@��t$@9w ~��O��� �E�L$@Qj ���$VPj�^� �����E�������ً] ��t�3����   ������A��   ���������Aug���������Au`���!��������AzS��~O�E �؅���]t��3ۃ  ~���3��O�'� �ESj ���$VPj� �E�����������ًE ��t�0�G��������Dz���E�D$D����ݜ$�   ݔ$�   ����؋] ����  ;t$H��  �O���ܜ$�   ����A��  ݄$�   �����A��  S���j��T$TR��$�   P�����$�����G��Sj��$�   Q��$�   R�����$�k����D$<����   ����   ��t��t	���  �L$L�T$P�D$T�L$d�L$X�T$h�T$\�D$l�D$`�L$p�L$|�T$t��$�   �D$x��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   �L$d��$�   ��$�   �X����$�   �X����$�   Q�L$h��R���](����zc�E$���D$+t�    �E����   �O����   �L$L�~V����4����$�   �$R��$�   P�L$\�9R������X����t�t$D�E�/����E�] ��u�D$<;�t4�E0�U$�E���\$���E(�$R�ESP���\$�$V�����D$+��؍L$,Ǆ$@  �����e� �D$+��$8  d�    Y_^[��]�0 ���������U������4SVW���O�D$;�� �����t$<��  �EP�=����W����E���щM������A�b  �������T  ������  ����  �E��t��3ۃ  ~���3��O��� �ESj ���$VPj�v� �O���D������� �������@� ��������4� ���@��������A��   �E�������!��������Az��~������]�f�a��������AzX�O�I� �N;�}I�W�E�D����]t��3ۃ  ~���3��O�� �ESj ���$VPj貗 ������؋]��t�3����   ;t$<}{�G���]����Dzk�MQ�I����E���E�����|N��~��	uD�]�E8��(�\$ �E0�\$�E(�\$�E �\$�E�$S���$Q���V����D$;_^[��]�8 �؊D$;_^[��]�8 ����������SUV��W�{��3��>� ����|m��������K������{3Ƀ�|;�V������G��    �@��� �����X��@����X��@����X��@����X�u�;�}�σ�;����\��|�   ������_^��][�������������SV��W�~2ۃ�|u�N�V����t;�F� �����\�����Dz"�F�@�\�����Dz�F�@�\�����D{.�F�L$�T$��L$�P�T$�H�L$ �P�T$$�H�P��������_^��[� ������������SW���G2ۃ�|V�4@�G����L0���U����t2�G� �\0�����Dz"�G�@�\0�����Dz�G�@�\0�����D{2�O�T$�D1�L$��T$�H�L$�P�T$ �H�L$$�P�H�^���<���_��[� ����U������tSVW���O3��X� ���D$�g  �M ��t��3�9w ~�O�3ɋu�ERV���$QPj�˔ ������؉\$t��ua�G�E�\$ �L$ �D���Q���\$� �$V�  ����t2�  �D$ �U~�G�3��T$SV���$PRj�`� ���D$�؋G�؍��T$0�@�T$(���E��������Dz
�����������������O�T$�[��ۍ4�FP���T$\�$R�M�����d$(��P�D$<PV���L$|�$Q��L������� L���D$8�u��   �D$@�^9W(u�D$H�^�M��|Z�G�UÍ4�P�T$l�HR�L���D$(�d$0P�����D$\�$P�L���D$`�M��D$h�   �^��9W(u�D$`�^��A����   |g�E���Y�����\$��   �\$ �\$���V9W(u�V���V9W(u�V���V9W(u�V���V9W(u�V��u��\$ ;�"�E��+�������V9W(u�V��u�E �؅�t�L$��   _^[��]� _��^[��]� ���������U����j�h]�d�    P��  SVW�  3�P��$�  d�    ��F �X����\$P��  ;F��  �}���B������  ��Ph��$�   Q���ҍ�$�   Ǆ$�      �fB�����H  ��O�W�D$T�G�L$X�T$\�D$`��$�   Q�L$XƄ$�  ��W�����L$T��  �B������  �T$T�D$X�L$\�T$<�T$`�D$@�L$D�T$Hj �L$XƄ$�  �D$8�����D$(�����@��� j�L$8Q�����$�H ��t*�D$4��|";��V��j �\$0�L$@�p@���D$,�j�L$X�_@��� j�L$(Q�����$�� ��t/�D$$��|';�#�V��j�\$0�L$@�!@���D$,��l$$�L$<�-A������  �L$4����  �D$$;���  ;���  ��������$�   P�L$@�]V����t}�~j �L$X�?��� ��N�4�j�L$X�?��� �L$<�Ƅ$�  �a� �L$TƄ$�   �P� ��$�   Ǆ$�  �����9� �   ��$�  d�    Y_^[��]� �S��\$$;�}�{W�N蕀��W�N茀�����\$P�|$4����  �D$P�^�N+ǃ�����$�   ��$�   �D$8    ���  �T�A0�эS�\���$�   �\$P+߃�������$�   �ۉ\$8ߋ�$�   �\$,��    �G��� �ZЋYЉXЋYԉXԋY؉X؋Y܉X܋Y��X��Y�X��G��Z؋Y�X�Y�X�Y��X��Y�X�Y��X��Y��X���Z����Y�X�Y�X�Y�X�Y�X�Y�X�G�Z�Y�X�Y�X�Y �X �Y$�X$�Y(�X(�Y,�X,��`�� ��`��$�   �A����|$4��$�   ��$�   �T$,;T$P^�D$8�@�<R�����|$8�<��|$8�Ӌ|$8�D$8��9�8�y�x�y�x�y�x�y�x�y�x������;T$P~��|$4�D$$+ǍxW�N�D$(�D$8    �~��W�N�~���F� j �L$@�\$0�,=��� �\$,����At'�|$$ u�~j�L$@���=��������At2����D$$;D$4~K�N����j�\$0�L$@��<��� �\$,����Au&�V�D$$j�L$@�|��<�����D$*����At�D$* ���-  �F�@���\$��$  � �$�VQ���F��L$d�P�T$h�H�L$l�P�T$p�H�L$t�P�T$x�H�L$|�P��$�   �H ��$�   �P$��$�   �H(��$�   �P,�D$|P�L$hQ��$  Ƅ$�  ��$�   �c� ��Fݜ$�   ��2��\$,j � �L$@ݜ$�   Ƅ$�  �\$/�;��� ܜ$�   ����A��   �~j �L$@���;��������Aukj �L$@�;��� ����$  �$��;��ݔ$�   ����$�   �$R��$  ��� ��L$d�P�T$h�H�L$l�P�T$p�H�L$t�P�T$x��|$$ ��   �F� j�L$@ݜ$�   �;��� ܜ$�   ����A��   �~j�L$@����:��������Auzj�L$@��:��� ����$  �$�;���T$,����$�   �$P��$  �5� ��L$|�P��$�   �H��$�   �P��$�   �H��$�   �P��$�   �D$+�D$,݄$�   ��������u}��$  ��Ƅ$�  ��� ��$�   Ƅ$�  �� �L$<Ƅ$�  �׈ �L$TƄ$�   �ƈ ��$�   Ǆ$�  ����诈 3���$�  d�    Y_^[��]� ����   ��4������   �D$|P�L$h�^X����;����Aze�|$$ ~^�F�@��j�\$0�L$@�r9��� �\$,����Au9�V�B�Nj �ЋV�B�Nj �ЋF�l$$� j �\$0�L$@�29���D$,��~j �L$@�9��� ��L$d�F��T$h�P�L$l�H�T$p�P�L$t�H�T$x�P��؀|$+ tT�~j�L$@����8��� ��F�L$|�H��$�   ���P��$�   �H��$�   �P��$�   �H��$�   �P��$  Ƅ$�  �K� ��$�   Ƅ$�  �7� �|$* �P  �L$$�F�D��ȃ��\$��$�   � �$�M���D$$�@�F�ЍЉ�$�   �P��$�   �H��$�   �P��$�   �H��$�   �P��$�   �H��$�   �P��$�   �H ��$�   �P$��$�   �H(��$�   �P,��$�   P��$�   Q��$D  Ƅ$�  ��$�   ��� j�L$@Ƅ$�  �z7��� ����$�   �$��7���T$,����$t  �$R��$H  ��� ��4��\$,��$�   �P��$�   �H��$�   �P��$�   �H��$�   �P����$�   ��ue��$�   P��$�   �U����;����AzD�|$$��~@�_S�N�'x��S�N�x���N���|$$�D��|��\$,j�L$@�6���D$,��|$$�Vj�L$@�|��6��� ��D$$�N��$�   �D@�����$�   �H��$�   �P��$�   �H��$�   �P��$�   �H��$<  Ƅ$�  ��� ��$�   Ƅ$�  �܄ �~j �L$X��5��� ��F �V�t���:��������������U����j�h��d�    P���   SVW�  3�P��$�   d�    �����   �҅�t2���$�   d�    Y_^[��]� �N�|� ��|ً]���6����tˋ�Ph�L$4Q���D$* ��P��Ǆ$      ��K���L$4�D$'Ǆ$   ������� �|$' t���$�   d�    Y_^[��]� �~j ���5���������   �F�@�D$&� �T$,���������3����FP��$�   Q�H��=���F��~�T$4�H�L$8�P�T$<�H�L$@�P�L$|Q�T$H�@j �ˉD$P�4���'����$�   �t$8�$R�7>����P�L$8��<���~j ���^4����L$4�F��T$8�P�L$<�H�T$@�P�L$D�H�T$H�P�N�� ���F����    ��L$(j�ˉD$0�4���D$,�����A�  �N�T$(�
�
�`��D$&�T$4�������������F�<�����Q�R�D$hP��<���F�8ǉL$L�P�T$P�H�L$T�P�T$X�H�L$\�P�FD$(�ˉD$,�D$dPj�T$h�h3���L$0�!����$�   �t$@�$R�=����P�L$P�;���FD$(j�ˉD$0�*3���D$,��F�L$L�8�T$PǉP�L$T�H�T$X�P�L$\�H�T$`�P��|$& t��蕶���D$&��$�   d�    Y_^[��]� ���������U����j�hɔd�    P��hSVW�  3�P�D$xd�    ��3��O�t$0�t� �؃�}�M�u���ƋL$xd�    Y_^[��]� ��P4SjV���ҋMP��t����t�3���~6�t$,�G���M���$V�i���OL$,Q�MV�f���D$,��;�|΋]��t2��Rh�D$4P����P��Ǆ$�       �D$4   ��G�����D$+u�D$+ �D$0Ǆ$�   ����t	�L$4�o� �|$+ �ut����   S���ҋ�Pj ���҅�t�   �L$xd�    Y_^[��]� 3��L$xd�    Y_^[��]� ��������VW�|$��t5h�X���
�����t%�t$��th�X��������tW������_�^�_2�^�������������j�h��d�    PQVW�  3�P�D$d�    ��t$肳��3��N�|$�L+�ޠ �F%�~�~ �~$�F(   �ƋL$d�    Y_^������j�h3�d�    PQSVW�  3�P�D$d�    ���|$�L+�w3�9^�D$   �%t�F;�tSP���%�^�^�^�O�\$�������D$���������L$d�    Y_^[���U����j�hv�d�    P��hSVW�  3�P�D$xd�    ���E�03�;��D$ �\$th�X��肔������   �t$�M�1��th�X���a�������   �ދG �p�����  �O�E�����A��  ��������  j�T$$R�����$���  �L$ ���D$}����  ����  ;���  �W�E�����A��  �������w  �|$ t �A�D$�3��L$xd�    Y_^[��]� �Q�T$�w �D$+�;���   ��u7j,�������D$��Ǆ$�       t	�������3�Ǆ$�   �����D$�D$�L$��P��s���L$Q�L$���o���T$�L$��R����D$�L$P���o���T$�G�L$�I���RPQ�S
 �D$$�P�D$(�O�@���PQR�4
 ���|$ t�L$���n����E��O(�T$�J(;���   ��u5j,�������D$��Ǆ$�      t	�������3�Ǆ$�   �����؍KV�s��V�K��n���KV�C��V�K��n���G �O+ƍ�    R��P�CP�	 �G�O�v�+�ҍ@�R���CQP�k	 ���|$ t�S�E��G(�C(�L$�E�A���\$�L$4� �$��A���L$�P���   Ǆ$�      �Ѓ���L$$��$�   �{ �K�O���� ���\$�L$D�E�$�A���P���   ��Ǆ$�      �ЍL$4��$�   �O{ �D$��؋L$�U�E�
��D$�L$xd�    Y_^[��]� ��������������U�l$��V��~Q�|$ tJ�FS�^W�<(;�~�n��;�}��;�}P�������T$�F��    Q�NR��R�+ ��n_[^]� ��������������j�h��d�    PQ�  3�P�D$d�    j,�������D$���D$    t�������L$d�    Y���3��L$d�    Y���������������j�hەd�    PQVW�  3�P�D$d�    ��j,�$������D$���D$    t���*������3����D$����t-;�t)W��輻���GP�N�u���V�R�N�GP�ҋG(�F(�ƋL$d�    Y_^����������V���8����D$t	V��������^� ��U����j�h)�d�    P���   SVW�  3�P��$�   d�    ���Ph�L$tQ���ҋ���   ��Ǆ$       �ҋ����|$L�"  �Ej ���T$`��$�   �$�~,����u=�E���L$|�$�h*�����k ��������Au��$���L$|�$�*���\$T�D$Tj����$�   �$�%,�����u  �N赢 �D$Tj j �؋F���$PSj�\$l�Ez ���F�����D$p����������z0�L$t��Ǆ$   �����2x 3���$�   d�    Y_^[��]� �Q����t��������Dz�\$H��K�L$H�T$HR��$�   �q���D$HP�L$hƄ$  �_����N��Ƅ$   �D$T��������Dz�F�؍�������$�   �$Q��� ����H���$�   �H��$�   �P��$�   ��$�   �P�@��$�   Q��$�   ��$�   ��$�   ����T$TR�L$h�Ss���F�L��+�R��S��$�   �Q���F�D�PS�L$l������D$H+D$P�\$l�|8��F��PW��$�   �`Q���F��PW�L$l������$�   Q��$�   ����T$TR�L$h��r���L$t�(��;\$l}�D$h�؃����\��;\$l|ꍄ$�   ��P�L$X��q���L$TQ�NƄ$  �0� �L$TƄ$   �����V�R�N�D$dP�ҍL$dƄ$   �n����$�   Ƅ$    �J�����D$L   �>�L$t��l�(���E������ɋ��\$�$�Ћ|$L�L$tǄ$   ������u �ǋ�$�   d�    Y_^[��]� �����������VW���T$���T$�$�.������T$�N�\$���$�.������T$��N0�\$�$�.������\$�NH���T$�$�i.���~`���O9�����Vx���Vh���_�^p^�������������D$��HV��W�F0P���L$�$Q�0���D$h�|$d��PW�VR���D$4�$P��/����P�L$DQ��� /������.����_^��H� ��������������̃��AHPQ�L$Q�L$(��.�����#/����� ������������̋QH���ĉ�QL�P�QP�P�QT�P�QX�P�Q\�P����ĉ�Q�P�Q�P�Q�P�Q�P�Q��`�P�7����������̍A������������̍A0������������̃�VW��V�D$P�L$,�J.���|$<��t�NQ�L$�e.����|$@��t��0V�L$�N.���_�^���  �̋D$��SUV����P�V�H�N�P�V�H�N�P�D$,�V��NH�P�VL�HW�~H�O�P�W�H�O�P�ωW�3���nW�͊��(������2��U�D$WP� 5����V0�P�N0�Q�P�Q�P�Q�P�Q�@���A��2�����{���_^]��[��� ��������������̃�S�\$$U�l$$�E V���M�N�U�V�E�F�M�D$0WP�N�US�~HU�ωV�B��U�L$Q�ˈD$4��,����V�H�n�M�P�U�H�M�P�U�@�͉E�2��U�L$WQ�A4����V0�P�N0�Q�P�Q�P�Q�P�Q�@���A��1����W���ĉ�O�P�W�H�O�P�W�H�P��V���ĉ�N�P�V�H�N�P�V�H�N`�P�=5����u
_^][��� �D$,_^][��� ̃�(SV��W�~`���5������   ��V���ĉ�N�P�V�H�N�P�V�H�ωP�6�����T$��;����AuJ����/�����Fx�����T$��'����Au ���]3����t�D$�h,�\$����z	2�_^[��(Í^H�F0SP��V�:?������tߋ�W�G�L$�O�T$ �W�D$$�G�L$(�L$�T$,�D$0�0���L$SQ�2���%�$������4����At�_^�[��(�����̃�SUV��n,�F�N�V �^(�l$ �n0W�~$�n�n4�n�n8�n �n<�n$�n@�n(�nD�F0�D$$�N4�V8�~<�L$�~HQ�^@�ωn,�FD�-�����H�O�P�W�H�O�P�W�@�ΉG����_^]�[��������V���H(���N�@(���N0�8(���NH�0(���N`��3���D$�L$PQ��������^� ̋D$��8SUV����P�V�H�N�P�V�H�N�P�D$L�V��N�P�V�HW�~�O�P�W�H�O�P�ωW�/���l$TWWU�1���$�D$$P�7*����P�L$4Q���)����V0�H�^0�K�P�S�H�K�P�S�@�ˉC�.��S�L$4WQ��0����VH�H�~H�O�P�W�H�O�P���W�@�ωG�~.���Ί��5�����t?��������؄�t2W���,)������\$�.����4�\$����z_^]2�[��8� _^]��[��8� ���������   VW��$�   ������$�p�����t������_^�Ĩ   � SV�D$@P���,����G`����������Dz<�Gh������Dz0�Gp������Dz&�Gx��$����Dz�NQ�T$XR�ϳ蒴���8�؍D$<P��$�   Q�VR�D$xP��2���'��P��$�   Q��诳������'����H�T$�P�L$�H�T$�P�@�ۉL$�T$�D$ [t�N0Q��$�   R�������1�D$8P�L$lQ�V0R��$�   P���h'��P�L$\Q���;������'����T$ �H�L$$�P�T$(�H�L$,�P�T$0�@�L$ Q�T$�D$8R�D$@P���5���_^�Ĩ   � ���������́�   SV��$�   2�����waW��$�   ��wSj�L$耭��V�L$薮����W���L$臮����V���L$�x�����W���L$�i��������ˍD$P�����_^[�Ā   � �����������́�   SV��W�L$$������$�   S����)��݄$�   �������8  ��=��=��$�   �� >�P�>�H�>�P�>�H��P�W���ĉ�O�P�W�H�O�P�W�H���P�\$݄$�   �L$d�$�l����sV�D$P�L$,�:������P�V�H�N�P�V�H�N�P�V�s0V�D$P�L$,�������P�V�H�N�P�V�H�N�P�V�sHV����(����u1V�D$P�L$,�Ʊ�����P�V�H�N�P�V�H�N�P�V���]���_^[�Ę   � ��V��N�P�V�H�N�P�V�H��$�   �P����ĉ�Q�P�Q�P�Q�P�Q�I�P�H���\$�L$d݄$�   �$�G����T$$R�������_^[�Ę   � ���������������V���"���N�"���N0�"���NH�"���N`�(.���D$�L$�T$PQR���R�����^� �����������̋D$�D$V��VP� ���$�D$�� �����$����^� ��������������j�hc�d�    PQVW�  3�P�D$d�    ��t$�D$   蚭���~��萭�����D$ 脭�����D$�����u����L$d�    Y_^������V���X����N�P���3��F�F�F�F�F�F�F �F$�F(�F,�F0�F4�F8�F<�F@�FD�FH�FL�FP^���̅�tf��t\�QV�p;�|A0�Q�p;�|5$�Q�p;�|)�Q�p;�|�Q�p;�|~�   ^Ë	� ;�}���^�3�;���^��ø   �����̃�$3�V��W�D$�D$�D$�D$�D$�D$�D$ �D$$�D$(�~,�ǍL$�D$   �D$F   �E������N���7�����_�   ^��$�_3�^��$�VW�|$j ��j���ͳ������tSV��讱������tD�FP���,�������t2�NQ��花������t �V,R����������t�FPP��趭����_^� �������������̃�VW���D����|$�D$P�L$Q���D$    �D$    �O�������tZ�|$uSV���I�������tD�VR����������t2�FP���%�������t �N,Q���Þ������t��PV��������_^��� ������j�h��d�    PQV�  3�P�D$d�    ��t$�D$    �۪�����D$�����̪���L$d�    Y^���������������˫����������̃�SUVW��蒪���|$,3ɉN�F�D$�N�F�D$�F��D$ �F��D$$�n�M �^��L$�L$�D$P�L$Q������������   �|$u|���)���S����������tfV����������tWU����������tH�T$R�����������t5�D$P���͚������t"�L$ Q��躚������t�T$$R��觚����_^][��� ����������VW�|$j ��j���=�������tw�FP���k�������teV����������tV�NQ���J�������tD�VR���8�������t2�FP���&�������t �NQ����������t�VR��������_^� ����������j�hÖd�    PQV�  3�P�D$d�    ��t$賩���N�D$    裩���N�D$薩���ƋL$d�    Y^������j�h��d�    PQSVW�  3�P�D$d�    ��t$�D$   蹨���~��诨���^��襨�����D$�I������D$ �=������D$�����.����L$d�    Y_^[�������������̃�VW�|$��D$P�L$Q���D$    �D$    贯������t/V��赝������t �VR��裝������t��V��葝����_^��� ������VW�|$j ��j���=�������t/V����������t �FP����������t��V���������_^� ��VW��������wT���=���3��Op�F�F�F�F�F�F�� ���   ���d����N�\���_�N^�R�����j�hL�d�    PQV�  3�P�D$d�    ��t$�D$   �{������   �D$�����Np�D$�� �NT�D$ �������D$����������L$d�    Y^���̋D$=���|�L$�A�h�,h�,h�  h|,��  �T$���B    �����̃�SVW��������t$�D$P�L$Q���N��������#  �I �D$=$�  wQt>-!�  t*��t����   V�Kp�� ��   V�KT�7����   V�������   V���   �����   =%�  ��   =&  ���   �L$�� �D$|=L�w���tP��L|=�L�sCh-h -h�  h|,��  ��3�h�,h�,h�  h|,��  ���F    �=���|ԉF�	V�Kp�N� ��������t.�|$�t�D$P�L$Q���+��������������_^[��� _^3�[��� ����������UVW��覗���|$Ph&  �����G�������G  �����������5  ���������t8j h!�  ���G�������  W���<����ϋ��C�����u
3�_��^]� ����   S�]T���b�����u2j h"�  ���@G��������   W���}����ϋ����������   ����   �Ep�P�]pj ���҅�t+j h%�  ����F������txW����� ����������t`��t^���   ���դ����u*j h$�  ���F������t8W��������ϋ��k�����t!��tj j����F������t���J�����u3�[_��^]� �����������j�h��d�    PQV�  3�P�D$d�    ��t$�����N�D$    �������D$�FP    �����ƋL$d�    Y^���������������́�4  �  3ĉ�$0  3�SVWP�ىD$�D$ �D$$�D$(�D$,�D$0�D$4�D$8�D$<�M( �D$�D$P�T$�( ����t�	   ���|$�{,�	   �t$h   �L$@j Q�� ���T$R�D$@P�D$�  �  ��uf�D$<�L$<�sQ���3����{P V���CP    让���{�	   �t$�CP�CP��$<  _^[3��� ��4  ��j�h̗d�    PQSVW�  3�P�D$d�    ���|$�a����wT3ۋΉ\$聢���^�^�^�^�^�^�Op�D$��� ���   �D$�r������D$�����ǋL$d�    Y_^[����2���������������V��3�9tc�h[��   ;�uV�5lc��2}:;�u�k4;�t8tRWQVhX.�^WQVh8.h�  hh[��� ���^Ã=hc2utVh�-�X��t��ub�5hc��2}:;�u�k4;�t#8tRWQVh�-h�  hh[�w� ���^�WQVh�-�uj2hh-h�  hh[�N� ���^��̸h[�P�����u�+�y2�ù�  +ȃ�|�T$R�T$RQ��h[P�gc �ޒ�������������̋hc�T$��2��=tc �hc�h[tK��2})��u�k4�D$PRQh�-h�  hh[�� ���uj2hh-h�  hh[�� �����t.�L$��t�9 t�T$RQ�&�������thh[j��| �����������������̋hc�T$��2��=tc �hc�h[ty��2}W��u�k4�D$��t&�8 t!P�D$PRQh�-h�  hh[��� ���;�D$PRQh�-h�  hh[��� ���uj2hh-h�  hh[�� �����t.�L$��t�9 t�T$RQ�H�������thh[j��{ ���̋lc�T$��2��=tc �lc�h[t��2}W��u�k4�D$��t&�8 t!P�D$PRQhX.h�  hh[�� ���A�D$PRQh8.h�  hh[��� ���!�=hc2uQh�-h�  hh[��� �����t.�L$��t�9 t�T$RQ�r�������thh[j �{ �������������̃|$ uQ�T$�L$�hcW�|$�   �K�����_t.�L$��t�9 t�D$PQ��������thh[j�z ���������̸�c�����������V���X����N8N$��8N ^���������̃y �At������3�9D$���D���|���� 3�� ���3�9D$���T��D�RP�XW ��� �̋A<��t�Q0�I4�T$�L$э�� 3�� �����������̋A<��t#�y t�Q0�T$V�q4�t$�Q^��� ��� �SV�t$��W��t�   �L� �\$;�}=�D�(��t��t1��    QP踻�������    R�F������D�(���#ÉD� 3�9D�(_^��[� ������V��N8W�|$;�}:�F<��t��t/��    QP�X��������    R�������F<���#ǉF83�9F<_��^� ���������̃�U�l$�E�F�M�N�~ �U�V�E�F�M�F�N�UW�Vt�����ȉF4�N0�}( tx�V�FRP��U �N ����;�}:�F(��t��t/��    QP褺�������    R�2������F(���#ǉF �F�NPQ�vU �N(��    �E(RPQ�1� ���}, tx�V�FRP�KU �N$����;�}:�F,��t��t/��    QP�&��������    R费�����F,���#ǉF$�F�NPQ��T �N,��    �E,RPQ�� ���}< ��   �V4�V�VR���C����~ �Ft���M4����D$�E0;F0�L$u.�F4;�u'�N���N�U<�F<���QRP�I� ��_]��Ë~<3�9F�D$~\S��l$ �]<��t�M0�ȍ��3�3�9n~-�T$RSW�� �F4�<ǋD$$��������;n|׋D$��;F�D$|�[_]���VW�|$��;�tW�.� W�������_��^� �������������́�   �  3ĉ�$�   S��$�   UV��F�N�VWP�FQ�N�nR�VPQRh�.S蹜���� 3��d$ 3������L��T�QR�jS PWh�.S荜���E�M �U���PQR���7���������|��~ ��<u��<P�F�FPh�<S�H������~< uhx<S�4������   h�   �L$j Q�� 3���9~~d���~h�&S������W�T$h|.R�D$ �� �F<����t�N0�ύ��3��N�T$R�VP�F4P�FQRP���E�����;~|���$�   _^][3��� �Ą   � ��QU��EW3�;ǉ|$#�L$;���  Php0Q�f�������_]Y� 9}<u%�L$;��f  PhP0Q�>����D$��_]Y� SV�t$�D$   �]�|$ �/  ����D$    }����   PWh0V�������   �K;�}����   PWQWh�/V�˚�����r�S��u��tgh�/V谚�����WVRQP��Z ����u��tCWh|/V苚�����2�S ������;�}��t ����PRWh8/V�a�������D$   �������%����|$ tX�}���E�Hu�ȋU�х��Xu�؋E�}0��;�|9U4}(;�|9]4}��t�E4PWh�.V�������D$    ^[�D$_]Y� ���������̋T$3�9D$��P�D$R�Q<P�A4R�Q0P�AR�QP�A�IRPQ��j ��(��� ��j�h��d�    P��4SUVW�  3�P�D$Hd�    ��\$X3�Uj���W�����;���  �FP��聗����;���   �NQ���k�����;���   �VR���U�����;���   �FP���?�����;�to�NQ���-�����;�t]�VR��������;�tKU��������;�t<U���������;�t-�L$�=P �D$P�ˉl$T�����L$���D$P�����P 9n(t�N�VQR�GO �����tU��視������t�F(PU��裖�����~, t�N�VQR�O �����3��tU���h�������t�F,PU���e������~ �Nt���~< �L$Xt#��~�V��~�F��~9N0|9N4|���3��txU����������tk��~g�~ �D$    ~Y��tU3�9~~:��t6�F<��t�V4�N0���L$э��3��T$XPR���ȕ����;~��|ƋL$��;N�L$|���ǋL$Hd�    Y_^][��@� ���j�h9�d�    PQVW�  3�P�D$d�    ���D$    �|$ ���D$    �P ���D$$���D$    �D$   t�   �T�(�OQ�L�WR�T�QR�V ���ǋL$d�    Y_^��� �U��������S�]�T$��VW����   �   9F��   9F��   �~< ��   �   +Í�3�98�D$~u������F<�\$t��t�N0�ύ����t�V4�׍��3��T�0�L$Q�NP�D�R�VPQR�H �D$0�D$(��������Au���T$��؋D$��;8|�_^[��]� �������������VW�|$����t	j ������|$��tj��������_�   ^� �������������̋D$��t�   �T�(R�T��D�RP�M ��� ��������̋D$��t�   �T$R�T�(R�T��D�RP�N ����� �U����j�hh�d�    P��hSVW�  3�P�D$xd�    ��}��PlW�L$8Q��3��ҍL$4��$�   �>���\$,�L$4����D$,������Azh3������L�(�T��D���t��E��������z���D����T������Au���D�����ʋE�ʋMPQ���\$���\$�$� �� ������؍L$4Ǆ$�   �����tL �ËL$xd�    Y_^[��]� �������������SUVW�|$4����t��3ɋl$0��t��t�   �����D$�VQ�NP�F(���$PQR��M ������t�O�3Ƀ�t��t�   �����D$�VQ�NP�F,���$PQR�M �D$8�T$H�N0��R�T$,R�T$,���\$���F4�D$,�$R�ы�����Ջn<�T� R�V(P�F,Q��Q�N�ڋVP�FQ�NRPQ�ax �L$t��@����t��y_^][�$ �������U����j�h��d�    P��   SVW�  3�P��$�   d�    ��}3ۅ�t	����  ��Pj �҅��t  �F3�9^t��j,�D$T�������D$T;É�$�   t!�L��T�Q�NR�VQR���Fk���؉\$L��\$L��Ǆ$�   �����X���K���P�D�(PQ��� �E��j �   +�j�   +Ǎ�������$�   +ωD$d� �<��RPQ�L �����D$D}
�D$D    ��T$T�
+;�~�L$D�?�L$LWWj ��� �D$\P�L$h�j���L$XǄ$�      ����T$t���P��\$H��QR�1� 3���9|$l�|$T��   W�L$\����M�|� �D$H    ��   �ɋN<t��t.�V4�T$H��~0������t�V0�T$H��~4����3ɋ\$P3���|2�S������<�    ��� �X��� ���A��X��A��X��A��X�u�;�}��+�����X�����u��T$H�M�\$D�|$T��;T��T$H�P�����;|$l�|$T�����t$L�F(j j P�L$d��r �EPj ���L$t�$�S*���L$XǄ$�   �����i���Ƌ�$�   d�    Y_^[��]� �Ë�$�   d�    Y_^[��]� �����������j�hۘd�    P��UVW�  3�P�D$$d�    �|$43���l$��  9k<��  �t$8;�u/j,�������D$ ;ŉl$,t	���:���3��D$,�����D$8��9k�kt���L��T��   +Ǎ��D$� ��QRj P���u;�����L  �N(;K<u�V �V���R�ª�����D$�F(�|� ��    �D$�D$    ��   �L$Q���>�����s<��t��t�S4�T$�4����t�C0�D$�4��3��L$3�99~>�   +T$4���D$ ��$    �L$QVU�d� �T$,�L$$�l$ ����;9�4�|ًD$�T$4�t$8��;D��D$���`����l$��t$�N �N�C<���QUP�F(�� U�������V;T�(t���N���N���P�D�(PQ��� ���ƋL$$d�    Y_^]�� �3��L$$d�    Y_^]�� ������������̋��{�����{����w	�W(3�;�u3��9Ou�9NU�nt���   +Ë���;Gt3�]�9N8~�F<;�t;�tP�T�����3ɋW$�V8�G(�F<�O$�O(9L� ~�D�(;�t;GtP�$�����3ɋW�T��G�D��W�T� �G�D�(�O�O�O �   +ӉL�0�,��   ]������j�h �d�    P��\SUVW�  3�P�D$pd�    ��$�   �   ;���   ��PlW�L$Q����j �L$�D$|    �1����5���$�   ����Dz5S�L$�����5�����Dz�E �M�U�D$�E�L$�T$�D$ �L$$�������RlW�D$8P�Έ�$�   ��PU�L$,Ƅ$�   �d���L$4�\$x�wD �L$$�������L$$u2�D$x�]D �L$�D$x�����LD 3��L$pd�    Y_^][��h� j �]���j �L$���P���� �] ����DzES�L$(�:���S�L$���.���� �] ����Dz#�L$$�D$x ��C �L$�D$x������C ��녋��x���L$D�o6���D$DPW��Ƅ$�   �Z�������t�L$$Q�L$H�uT����t�ߍ|$D�V����L$D�D$x�d���L$$�D$x �jC �L$�D$x�����YC �   �������������������j�hH�d�    P��0SVW�  3�P�D$@d�    ��|$P3ۃ��\$��   ����   W�҅�uv�L$�5���D$P�\$LW����������t+�L$TQ�L$��W���ߍ|$�D$�����|$ t���w���L$�D$H������c���D$�L$@d�    Y_^[��<� 2��L$@d�    Y_^[��<� ���������V�t$Q��������   ^� ��������̃�SVW�|$$�����D$ ��   �~ ��   �D�(�L��T�jPQR��F ��������   �F<U�nj ���U�D$�3����^3Ʌ������S�D�j �������������S��U�ΉD�������L$�V�؋D$P�FQRP�V ����]tU�L$�V�FSQRP�; ����t;�N<�V4�F0WQ�NR�VP�FQ�NRPQ�# �� �����   W�Ѕ�t�D$�D$_^[��� ����������̃�S�\$��UVW���D$ wI�D�(�L��T�PQR��D �����D$t*�D��|����   +ˉD$3�����9�D$�L$�D$_^][��� ��\$$�ۋn<t4��t,�V0�N4����э\� ��tN�V0�N4���L$эl� �:3����t,�V4�N0����э\� ��t�V4�N0���L$эl� �3���3��|?��$    �V�FUSRP�� ����tD�L$$�D�0�l$�����+�+��}̋D$�T$��;�D$�5����D$_^][��� _^]3�[��� ����������UVW���t���F<���   t�N0�V4�L$�T$ʍ<ȅ�u_^3�]� �D$������  �$���
�F�L$���PQW��� ���~ tk�V���׋�_^]� �~ �T$t�F��   QRW�� ��_^��]� ��S�^��������D{�4�3Ʌ�[~��+����Ƀ��X�;N|���_^��]� �~ �T$t0�F��3Ʌ�~��+����Ƀ��X�;N|�F��_^��]� �N���QRW�� ��_^��]� �~ �vt��L$��    PQW��� ��_^��]� _3�^��]� ��
��
_�
��
��������V���(s���N<3���tN�V0�T$W�~4�|$׍х�_t3�D$� ��~~�@�Y�~~�@�Y�~ t��F���   ^� �������������VW���r���F<3�����   �N0�L$�V4�T$ʍȅ���   9~t3�D$� ��~~�@�Y�~~�@�Y�V�@_�Ѹ   ^� ��T$�Z������D{�r�   �����~~"�B�����Y�~~�J_^�Y� _��^� �؋�_^� ���̋A<V3�����   �Q0�T$W�y4�|$׍Ѕ�_��   9qtX�A��������D{z�A���4D$�����y~�B������X�y~��^�J�X�   � ��^�X�   � ��D$��y��~�B����X�y~���B�X�   ^� �؋�^� ��������������D$<�D$�T$��(�\$ �D$\�\$�D$T�\$�D$L�\$�D$D�$P�D$<���\$�D$D�$R襮 �@ ��VW�|$����wSS��p���D�(�L��T�PQR�C �N4�V0W�؋F<P�FQ�NR�VPQRj�& ��,��[t��t
_�   ^� _3�^� ���������V���hp���F�N�V�F�F�F�F0�N�N4�F4�F �V�V$�F$�F(�N0�N,�F,�V �N(�   ^������QSUVW���p���F�N�   3�;��T$W����   �\$�l$�F<��t�N0�ύ��3��V4SUP�FRP� ����u�D$    ��;~|ŋD$_^][Y� ��~O�\$�l$�F<��t�N4�ύ��3��V0SUP�FRP�� ����u�D$    ��;~|ŋD$_^][Y� _^]��[Y� �����������j�hx�d�    P�� V�  3�P�D$(d�    ��~ ��   �o���L$�r� �N�F�V�L$�N0�D$�F�L$�N8�T$�V4�D$�F<�L$$�L$�D$0    �T$�D$ �� �T$�L$�D$�V�T$ �N4�L$�F0�V<�D$     �D$0������ �~ ���L$(d�    Y^��,������������̋�� �0����������0����������U����j�h��d�    P��hSVW�  3�P�D$xd�    �����Ph�L$4Q���ҋ�Ph�L$$Q��Ǆ$�       �ҍL$4Ƅ$�   ������\$�L$$������\$j����Az/�>�L$8�����j �L$8�����������\$��� �Gl�$���-�7�L$(�����j �L$(��������Vl���\$��� �$�҅��L$$��Ƅ$�    �\8 �L$4Ǆ$�   �����H8 �ËL$xd�    Y_^[��]����U����j�hؙd�    P��   SVW�  3�P��$�   d�    ���ڋC;G~����   ���Ћ������   �Ћ�P�]���K;O��  �ϋ��k�������  �s�L$t�t$P�������Ǆ$�       �a���ωD$L�V���L$L�D$T�6+T��T$X���   ���҅�u����   ���҅��R  ���3Ʌ��D$K~&�|$K t�W�C��������D{�D$K ��;�|ڋK�D$L�w+�����   ;t$T��   �|$K ��   �G�ȋS������D{�D$K ��;t$T��   �|$K ��   �G�D��\�����D{�D$K ��;t$T��   �|$K ��   �G�D��\�����D{�D$K ��;t$T}j�|$K tj�G�D��\�����D{�D$K �T$L�������;��9���;L$L}1;t$T}+�|$K t+�W�C��������D{�D$K ����;L$L|π|$K uJ�t$Pj���"(����tj���(����u0�L$tǄ$�   ������5 2���$�   d�    Y_^[��]Ët$P����S���;�|�G��;���  �G�D���K�\������D��  ;���  �W��;���  �������T$d�@�������D�j����W����T$l�@�������D�M����CVQP�D$\P��3 �O�WVQ�D$d�D$hRP�3 ݄$�   ݄$�   �D$t�у� ������   �O���؍�� ���\$��$�   �@��$������W��L$t�D$\�����D$\�@�j��L$x��� ������4�\$`����� �d$\�D$d��������u>�L$T�;��}�W��;�|��؋G���WV�\$pP�D$XRP��2 �D$d��   �D$X��P������D$d�L$LQ�����$�A���������A��   �K�����\$��$�   �@��$������S��L$t�D$\������D$\�@�j��L$x��� ������4�\$`������ �d$\�D$l����������   �L$L�;��}�S��;�|��؋C���SV�\$hP�D$XRP�2 �D$\���D$l�\$d����D�]����D$L�L$T;�~b�L$XQ������D$d�T$TR�����$�@�����'����D$T�D$L��K����D$X��P���k���D$l�L$TQ�����$�u@���^���}*�L$XQ���B���D$d�T$LR�����$�L@���������t$L������C;G��������X����3Ʌ�~"��[+���;����D���������;�|�L$tǄ$�   �����J2 ���$�   d�    Y_^[��]���j�h�d�    P��XSUVW�  3�P�D$ld�    ����f���L$�$��3ۍL$@�\$t�$���F<;��D$tt	9^8u�D$<�F(;�t	9^ u�D$0��$�   ��L$|����   R���T$ �$R��;ÉD$|%�L$@�\$t�R���L$�D$t�����R��3��(  ��$�   �$�   ����   P���D$L�$P��;É�$�   �L$@~��T$������t��D$(;D$Tu��L$$;L$Pu��L$�   �A[ ;�~�L$�4[ ���L$@�)[ ;�~�L$@�[ ���L$�[ ;�}�L$��L$@��Z ;�}
�L$@W�p ���L$�G�����L$@u�:����t	�L$���3�9\$ ��;�t	�D$�\$ �D$� Q�L$�$ ���F<;É|$�l$ t9^8~	P�ړ�����D$8�T$<�F8�F(;ÉV<�\$8t9^ ~	P賓�����L$0�T$,�   U�N(j�ΉV �\$4������F,��N,���Y�D$$�T$ �L$(�F�D$4�F0�V�+~��3�;ˉn�N�n�F4~OW�L$D����΋��d���F<;�t-�N0��N4��;�t9^�Ft����    RUQ��� ����;~|��t$|��$�   ;����L$@�\$t�P���L$�D$t�����P���ƋL$ld�    Y_^][��d� �������V�t$��th�c���+E����t��^�3�^����������������VW�|$��tBh�c����D����t2�t$��t*h�c����D����t;�tW��袔 W�<�����_�^�_2�^����������������V����~ ��0�xc3�;�t��F�F�F�F�F�F�F �F$�F(�F,�F0�F4�F8�F<��^�������Q�D$SUV��W�^SjP��� �NQjP��� �NQjP��� �~WjP��� �?��0������   �F���}   �~0 ~w�~4 ~q�~< tk�~ �t����    �L$3Ʌ��L$~K�~<��t�V0�э<��3�3ۅ�~%�D$WPU�c� �N4��F����;؍<�|ߋL$��;N�L$|��V�FRP�, �N(Q��    RU�� �N���FPQ��+ �V,��R�PW��� ��(_^][Y� ���̃� SVW�|$0��L�2ۃ�|T�T�;�|L�F(��tE�D$<�D$4������z0�D�(�D���T$�D���T$��������Dz!��������Dz���������_^��[�� � ������Au���W������������\$ ����$�\$(�����D$4���D$<3Ƀ��D$�D$�D$�D$$��   �Z��D�(�������D�(�ȍ�u���������������D�(�T������D�(�D��D�u���������������D�(�T������D�(�D��D�u���������������D�(�T������D�(�D��D�u������������Ń��;��L���;�}/�D�(�������D�(�ȍ�u������������Ń��;�|��ً��ڳ���������X`��_^��[�� � ������������V���8`���D$��}3�^� U�l$��}]3�^� W�|$��}_]3�^� S�\$$;�|�T$(;�}	[_]3�^� 3�9L$�F���n�~�^�V�ɉNt���F4�F0��P��Q�f) ��Pj ���i����V���FRP�J) ��Pj���M�����u3��N4�N�NQ��������u3�[��_]^� ����̋A<SV3�;�Wt	9q8t���3ҋA(;�t	9q t���3ۋA,;�t	9q$t���3�;։q�q�q�q�q�q�q �q$�q(�q,�q0�q4�q8�q<t	R聍����;�t	S�t�����;�t	W�g�����_^[�VW����^���|$W���>���~ u+���W`����Dz�Wh����Dz�_p����D{��؋��J����F<�N4�V0WP�FQ�NR�VP�FQRP� �� _^� j�h8�d�    P��`SUVW�  3�P�D$td�    ���2^����$�   �D$8P�L$ 3�Q�͉\$$�\$@�u����;���  �|$�z  �T$4R�͉\$8�\$4�\$0�\$,�\$(�\$$�\$@�\$D��]����;���   �D$0P����]����;���   �L$,Q����]����;���   �T$(R���]����;�t|�D$$P���]����;�ti�L$ Q���]����;�tV�T$<R���p]����;�tC�D$@P���]]����;�t0�L$D�' �L$DQ�͉�$�   �*^���L$D���D$|�����( �T$ �D$$�L$(R�T$0P�D$8Q�L$@RPQ������;�$�   tB��$�   R����\����;�t,��$�   PS���p�����;�t�O(��$�   QR����\����;�$�   tC��$�   P���\����;�t-��$�   Qj���"�����;�t�W,��$�   RP���y\����;�$�   t��$�   Q���L\����9_t�_���\$�	�W�T$�څ�t����$�   P���)�������$�    ~k��~g��ti� �D$    ~U��tW3�9_~:��t6�G<��t�O4�W0���T$ʍ��3�P�D$P����[����;_��|ƋD$��;G�D$|�3�;�u�������ƋL$td�    Y_^][��l� �������������j�h��d�    P��   SUVW�  3�P��$�   d�    �鋼$�   ���4  �E �PlW��$�   Q����݄$�   j��3��$�ȉ�$�   ��������$�   ��Ǆ$�   ������% ����   ��$�   � ���t$�t$t P���������D$��   ���Z���t$��$�   ���tP�S��������D$��   ���]Z���L$|����L$PǄ$�      � ���L$$Ƅ$�   �����T$|RW��Ƅ$�   ����������L$$uPƄ$�   �BF���L$PƄ$�   �1F���L$|Ǆ$�   �����F��3���$�   d�    Y_^][�İ   � ݄$�   �D$P�T$ �D$R�D$ P�L$(����$�   �$�<������   ��u3j@�m�����D$��Ƅ$�   t	��������3�Ƅ$�   �D$��;�t|�M�N�U�   +����V�(�0�   +����(�   +�S�͉0�P���PS��������   +�$�   S�����/����7���P�/PQ�[� ��$�   ���ߍ|$P������u7�L$;�t!��$�   ;
t��t��Pj�ҍL$$�����4����L$$�|����t$��u3j@�l�����D$��Ƅ$�   t	��������3�Ƅ$�   �D$��;�t|�E�F�M�N��$�   �   +����(�0�   +����(�   +�S�͉0�H���PS�������   +�$�   S�����'����7���P�/PQ�S� ����$�   �|$$������u\�L$;�t��$�   ;
t��t��Pj����5����L$;��������$�   ;��������������Bj�ЍL$$�Q�����$�   �8 u�L$���$�   �8 u�T$��L$$Ƅ$�   �kC���L$PƄ$�   �ZC���L$|Ǆ$�   �����FC���   �!���������������j�hۚd�    P��0  SUVW�  3�P��$D  d�    ��L$����3ۍ�$�   ��$L  ������$  ������$�   �������$�   �������$�   �������PlS��$�   Q���ҋ�Plj��$  Q��Ƅ$T  ����$SS��$�   P��$�   Q��$�   R��$�   P����$$  �$Ƅ$l  �d������\$��$  ��$�$�H��������$苀 ��;�t ��$�   �Y�����D����z3���  ��$�   ��$�   ��$�   �L$��$�   �T$��$�   �D$��$�   �L$ ��$�   �T$$��$�   �D$(��$�   �L$\��$�   �T$`��$�   �D$d��$�   �L$h��$�   �T$l�D$p���������   ��$�   ��$�   ��$�   �L$,��$�   �T$0��$�   �D$4��$�   �L$8�L$,�T$<Q�T$`�D$DR��$4  P�������L$P�P�T$T�H�L$X�P�T$\�H�L$`�P���L$D�T$X�_����L$������   ��$�   �E�������   ��$�   ��$�   ��$�   �D$D��$�   �L$H��$�   �T$L��$�   �D$P�D$\�L$TP�L$H�T$\Q��$4  R������L$8�P�T$<�H�L$@�P�T$D�H�L$H�P���L$,�T$@�����L$�f������$�   P��$�   Q�L$�����D$\������;�����D$l������4u_�D$d��������AzP��������������Az?�����������T$<�T$T�T$\�T$d��������Au���0'�L$�\$l�Ω����   �D$d��������AzZ����������AzM������������Az>�������������T$,�T$D�T$d�T$l��������Au���0'�L$�\$\�b����q������������AzR����������AzO��������������AzB���T$4�T$L�T$l�T$\�\$d����Au���0'�L$�\$d��������������������9^~S��ti3�9~~@��t<��$  RWS���:�����$  P�L$艨����ܜ$X  ����Au3��;~|���;^|���t��$T  ��t�    �t$󥍌$  Ƅ$L  �� ��$�   Ƅ$L   �� �L$Ǆ$L  ������ �ŋ�$D  d�    Y_^][��<  � ���U����j�h�d�    P��h  SVW�  3�P��$x  d�    ��3���$�   ��$�   �����L$<�n�����$�  ��$$  �   ����������y�$�  �   ���y�������y�$�   �e�����$�   �Y����L$\�P����L$t�G����}������<  �L$L�����l  ���  ���  �D$8�E$�L$T3�;��T$Xu��$�   ��$�   ��$�   �E$�](;�u
��$�   �](�U ;�u
��$�   �U �M���i  ��u3�E4���\$�E,�$S�EPR���\$�E�$QW���)� ���T	  �E�]����D�   �|�Q�4Z������Q�L$0�Y���ȃ����M�&  ���  ���  �D$% ���D$& �D$' u�D$'�D�3�8T$%�D$P   ��+Ѓ��T$4u�D$4    �M$�E��L�(R�T�j���$QRP�M �T�(���D��\�����ʍ�������\��@� ������4�E�E�������e  �T�����zw�D�������zj�D�����������Az[�T��C;�}P�M$�ً	�؋D�(�D�Qj�U���$P�D�RP� �E�E��������D$%������D$&������ڋU$�
�D��T��L����;ʉL$ }.�D�(������������u
����;�|�;��ɉL$ ��  �M9L$,t\�D��T�(�D���L��������AuC�����u:�E4�E(�M$�U ���\$�E,�$P�D$@QR���\$���$PW��~ ���'  ���؍L$<Ǆ$�  ������ 2���$x  d�    Y_^[��]�4 ������Au^��������AuR���$���������AzD�D����;�~9�M$�ً��؋��R�Uj���$P�D�P�D�P�H �E�E������ڋU$�
�D��L��P�;ʉL$ }(�D�(������������Az
����;�|�L$ ��;�k�M9L$,�����D�(�Ѝ�����������������������E4�M(�U$�E ���\$�E,�$Q�L$@RP���\$�$QW���} ����  �T$4���D$P�����T$4�D�(�����D$0�L$(����Au=�\$P�L$ ��~v�D��X�;�}&�T�(T$(�B�����Dz
����;�|�;ˉL$ |v�D$,2�;E�`  �E4�U(�M$���\$�E,�$R�U QR���\$���$PW�} ���.  �D��X�;�~��T�(T$(�B������Dz
����;��;ˉL$ ~��L$ �D�(�T$4���������D�4  �}�����V  W��$�   �����T$0�L$ �ʹ   ��   +ǋ�+ϋ�������;��D$(    �\$0��$�   ��  �   +Ǎ���$�   �	��$    ����$�   ��D��؃��\$�L$L� �$�����D$(���D$(�U  3ɸ   +�8L$%��$�   ������$�   ���$    ��$�   R��$�   ������D$(���L$D��$���$������M$���$�   ݄$�   ����   Qj��$,  RjS���\$��݄$�   �$�ЋE$݄$�   ����   Pj��$�  QjS���\$��݄$�   �$�Ҁ|$' ��  �\$&��tC�T$X�D$\P�D$P��$�   QRP�� �D$d��$�   Q�L$L��$�   RPQ�� �� �   �D$L��H��$�   �P��$�   �H��$�   �P�@��$�   ��$�   �D$8���$�   �P��$�   �H��$�   �P��$�   �H��$�   �P��$�   ��$�   ��$�   ������$�   ������$�   P��$�   �����E,��������A�  ���U  �E4�L$t�T$x��(�\$ �ă��}�\$0���$�   �P��$�   �H��$�   �P��$�   �H��$�   �P��$�   �ĉ��$�   �P��$�   �H��$�   �P��$�   �H�Pu�T����=����@����   �U(�L$ �   �D�(�ȋU ��!  �\$L���������4�D$8���$P��$   Q���������������2  �|$% tV�\$X��������4�T$T���$R��$  P���H������������u �M(�D$ �   �T�(�M ��   �؋D$(�����D$(������\$0��$�   �����;��D$(   �\$0�R����E�L$ �E�\$P�T�(ˍ�    ��D$(�L$ �T$0����A����������E(�    �T�(�ʋE ��L$<Ǆ$�  ����� ���$x  d�    Y_^[��]�4 �M(�؋D$ �   �T�(�M �뵋E(�T$ �    �L�(������؍L$<Ǆ$�  ����� �Ë�$x  d�    Y_^[��]�4 �D$��V����   �$���
�F,�N�Vj PQR�6 ��������t$j j ��诸���N�V0P�FR�VQRP�I� ����^� �F(�N�VjPQR�� ��������tڋFj ��P���`����N�V4믋N,�V�FjQRP� ��������t��N��Q�u����V(�F�Nj RPQ� ���������t���j j ��������N�V4�K���2���^� �I ��
�
8�
c�
���������D$V����0t	V�[������^� �U������tSVW���=E���]��P4���ҋu�D$X��P4���ҋM�D$\��P�ҋM�D$d��P��;D$X~'h2h�1h�	  h�0趴����3�_^[��]� �M��P��;D$\~'h�1h�1h�	  h�0������3�_^[��]� ���:������ΉD$T�,����|$T ���D$lu���D$L    t�D$L   ���C� �ΉD$P�8� �L$PPQ�ΉD$p����P�������T$XP�D$tRP��������O(;Kt%�W�GRP�� �S��    �G(QRP胜 ���O,;Nt%�W�GRP� �V��    �G,QRP�V� ���|$P �D$H    �m  ��]�L$HQ������3�9\$h�D$`�7  S�������ȋG<��t�W4�w0���t$H֍4��3��|$T t�D$X�T$`���T$x���
�����T$x�Ƀ|$l t�D$\���T$p����������Dz��������T$p����������������Dz�����������E��RVQ�L$h���$Q�����$�҄�������|$L tc�T$d�D$p�L$x3Ƀ�|7�B�������    ��� �����^����N��^����N��^����N��^�u�;�}��+���������^�u���u��;\$h������D$H��;D$P�D$H�����_^�   [��]� �����j�h;�d�    PQ�  3�P�D$d�    j@�HV�����D$���D$    t���n����L$d�    Y���3��L$d�    Y���������������j�hk�d�    PQVW�  3�P�D$d�    ��j@��U�����D$���D$    t����������3����D$����t;�tW���\r W��������ƋL$d�    Y_^������������������j�h��d�    PQ�  3�P�D$d�    j@�HU�����D$���D$    t���n����L$d�    Y���3��L$d�    Y���������������j�hțd�    PQV�  3�P�D$d�    ��t$�\ 3���0�xc;ȉD$t��L$,�T$(�F�F�F�F�F�F�F �F$�F(�F,�F0�F4�F8�F<�D$0P�D$(Q�L$(R�T$(PQR��������ƋL$d�    Y^��� �������V����0������^�[ ����������V����0�������[ �D$t	V�V������^� �����V�t$��thpd���� ����t��^�3�^���������������̸pd�����������VW�|$W���r���~ t�N��P0W�҃~ t�N��P0W�ҍN(�x
 _^� ���j�h��d�    PQV�  3�P�D$d�    ��t$�Z ����T$�T$�N�$�D$,    ��2�-����N(�e	 �hd��t��F    �F    �ƋL$d�    Y^������������SVW����P0j�ҍw�   ���t��Pj���    ����u�O(�	 ����T$�T$�O�$����_^[����������VW���=���~ ��t�N��P����~ t�N��P�����_^�������������V��~ t�N��T$�@R����D$�~ t�N�^�D$�B��^� ���������QUV�t$��;���   SW�����ݍ~+��D$   �? t*���Pd�ҋ�V�c<�������;u��t��Pj���҃��l$uǋD$�H�M�P�U�H�M�P�U�H �M �P$�p(�}(�   �U$�_[^��]Y� �S�\$UV��W3��u��> tN���P4�҃�u\���PS�҅�tv������|ԍM�<�����u{��th�3S��O����_^]3�[� ��tWh�3S�O����_^]3�[� ��t�L���P4��PWh�3S�O����_^]3�[� ��t�Whh3S�iO����_^]3�[� _^]�   [� �SV�t$WV���������N��h@4V�/O�����CP����R��h�&V�O����3����; Wt(h04V��N�������sN�����BV�Ћ��N���h4V��N����������|�_^[� �VW�|$j ��j���R������t=�FP���N���N(Q��� q������t �VR���>�������t�FP���,�����_^� ���̃�SUW�������\$�D$P�L$3�Q�ˉl$�l$�TR����;���   �|$��   V�WR���2<����;�t�G(P���0<����;��l$t7�L$Q���I����;�t%�T$R�9����;ŉGu�L$;�t	��Pj��;��l$t7�D$P���
����;�t%�L$Q�z9����;ŉGu�L$;�t	��Bj�Ћ�^_][��� ���V��3�9Ft,9Ft'�N��P4W�ҋ���~�N��P4��;�t_3�^Ë�_^��������̃�(�h ��������U����j�h>�d�    P��   SVW�  3�P��$�   d�    �ٍs(������������D$�h  �L$L�Z �L$|Ǆ$�       �F �K��Ƅ$�   t �D$P�o ��   �|$L�L$� �K��t �T$R��n ��   �|$|�L$� �L$L�G�������   �L$|�6�������   �sV��$�   P��$�   Q�T$(R�L$\�|������u�����K(�P�S,�H�K0�P�S4�H�K8�PV�D$ P��$�   �S<Q��$�   R�L$t�3������,�����K@�P�SD�H�KH�P�SL�H�KP�P�ST�s(���������L$|�|$Ƅ$�    � �L$LǄ$�   ����� ���*  ��P4���ҍL$�D$�� �} Ǆ$�      t\�E��tU�}��tN3�+ǉD$;t$},V�L$ �^����L$�9V�L$8��K�����������|΍L$���������   �s(�   �|$��B4���ЋU�]�ȋ�3�+ÉL$���D$;�};��tV�L$ ������ �L$���tV�L$8������ ��L$�U������|���~#��C�����t�t$�0��t�����u��؍L$Ǆ$�   �����q �D$��$�   d�    Y_^[��]� �C(P�L$ � �6������V��~ �t�N��PH�҄�t�~ t�N��PH^��^�����SV��~ �t(�N��PH�҄�u��P0j���ҋN��PL�҄��Ã~ t5�N��PH�҄�u'��P0j���҄�t�N��PL�҄�t^�[�^2�[�^��[������������́�  SV���P0Wj�ҋ�$  W���-���L$$3��¹���L$蹹���L$<谹���N��t@�D$TP�/I����L$$�P�T$(�H�L$,�P�T$0�H�L$4�P�N�T$8��PDW�ҋ؋N��tB�D$TP��H����L$�P�T$�H�L$�P�T$�H�L$�P�N�T$ ��PDW�҅�u3��   ����   U�nU�L$D�����D$P�L$\Q���F��P��$�   R�D$0P��$  Q���F��P��$�   R�D$PP��$�   Q�T$(R��$�   P�L$H�y������r���P��$�   Q���BF����苺����脺��P���\���]�~(���!  �T$lR���Ej ��   �L$l���  _^��[��  � ������D$V�D$����2�����z@�D$��w7�|� t0�L��ɋ�PlS���\$�$�҅���P0j��������[^� ������^� ���������������j�hy�d�    P��VW�  3�P�D$ d�    ���D$    �t$0���D$(    �N����D$4���D$(    �D$   u
9Gt>�O���u4� t.�O��@h�T$R�Ћ��P�V�H�N�P�L$�V���  �ƋL$ d�    Y_^�� � �������������U����j�h��d�    P��   SVW�  3�P��$�   d�    �E��U3��D$,   �D$<�T$@3ۍy�D�<;��6  �97u�t$,��\$4�t$0��@h�T$DR�Ћ���������L$T����T$X����D$\����L$`�L$l��$�   �T$d�D$h�I����t$(��I �D$(�L$0Qj ����T$tR���L$X�$��������$�8����t[h���L$X�L�����t�D$lP�L$X�z����D$4�\$4�L$l�T$p�D$t�L$T�L$x�T$X�T$|�D$\��$�   �L$`�T$d�D$h����@�t$(�_����D�<�D$4�L$D�Ǆ$�   �����!�  ��3�������������؋D$,��$�   d�    Y_^[��]� �T$3���u9At!�I��Px��� ��u9At
�I��Px��� ������������̋T$3���u9At+�I��T$�@|R��� ��u9At�I��D$�R|P��� ��̋T$3���u9At'�I����   ��� ��u9At�I����   ��� ������̋T$3���u)9AtO�T$�D$�I����   R�T$R���$��� ��u&9At!�D$�D$�I����   P�D$P���$��� ���������������U����j�h�d�    P��h  SVW�  3�P��$x  d�    �ٍL$D�Ӆ��3��L$,��$�  �ѳ����$�   �ų����$�   蹳����$�   譳����PlV��$  Q���ҋ�Plj��$   Q��Ƅ$�  ����$VV��$�   P��$�   Q��$  R�D$@P����$<  �$Ƅ$�  �1������\$��$4  ��$�$���������$�XZ ;ƉD$(�   ��$�   � ����%�$���p&����Au	�t$(��  �L$,�T$0�D$4�L$D�L$8�T$H�T$<�D$L�D$@�L$P��$�   �T$T��$�   �D$X��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   貹������   ��$�   ��$�   ��$�   �L$\��$   �T$`��$  �D$d��$  �L$h�L$\�T$lQ��$�   �D$tR��$4  P�~������$�   �P��$�   �H��$�   �P��$�   �H��$�   �P���L$t��$�   �����L$D辄����   ��$�   ��������   ��$�   ��$�   ��$�   �D$t��$�   �L$x��$�   �T$|��$�   ��$�   ��$�   ��$�   P�L$x��$�   Q��$4  R谺����L$h�P�T$l�H�L$p�P�T$t�H�L$x�P���L$\�T$p�K����L$D�������$�   P�L$0Q�L$L躄���};�t�    �t$D�3��s�I �|$( ��   ���$,  R�&@����L$D�P�T$H�H�L$L�P�T$P�H�L$T�P�L$D�T$X脃���E�����   ���T$L�$R�Ѓ������D$(|���tK�}��tD�L$,�T$0�D$4�L$D�L$8�T$H�T$<�D$L�D$@�L$P�L$D�T$T�D$X�����    �t$D󥍌$  Ƅ$�  �x�  ��$  Ƅ$�   �d�  �L$DǄ$�  �����P�  �D$(��$x  d�    Y_^[��]� ���̋T$3���u9At'�I����   ��� ��u9At�I����   ��� ������̋T$3���u9At'�I����   ��� ��u9At�I����   ��� �������3�� ����������̋T$2���t��uZ�|� tS�D$ ��t���3��D$0�L�����   V�t$(���\$�D$<�$V�D$,P�D$8P�D$(���\$�D$<�$P��^�4 ����U������4SV��3�9NW���   9N��   �];ىL$8�L$<t��K%��  �D$8�L$<�E@�N��}���   ��(�\$ �D$`�E8�\$�E0�\$�E(�\$�E �$P�E���$W�҄�tA�E@�N����   ��(�\$ �T$d�E8�\$�E0�\$�E(�\$�E �$R�E���$W�Ѕ�t�L$<�T$8������  ʉ_^[��]�@ ��������������̋D$VW3�����u
9~t�N���u9~t�N����   �ҋ�����)����_^� ̋A�Q�Q�A��)���   ����������U������4SVW����P4�|$03��ҋ�;��-  �E(;É\$8�\$<t��P����  �L$8�T$<�]���ދ���P�W���؉D$(�E$��������L$ w(�$������D$   ������   �D$�����	�   �D$�O�E�}(����   ����\$8#��]WP�D$,PVS���$�ҋ����G  �E(�E�|$0����L$<#��O����   P�D$ P�D$(PVS���$�҅��D$0�  ���] �D$    ~P�D$$���|$,�|$ ��+��D$(��+��D$4�D$�L$,P�e����L$(�9�D$�T$4�����;ƉD$�\:�|Ϻ   9U�T$,��  �҉T$(�D$    �n  �E���؅�~�΁�����3�������   �|$ �$  3Ƀ�|U�L$$�֍~������эC��    ��    ��� �@��� ���X��B��@��X��B��@��X��B��@��X�uҋT$(;���   �|$$����������    � ���D����;��\��|��   �|$����   3Ƀ�|V�L$ �����~������C��    ��$    ��� �@��� ���X��B��@��X��B��@��X��B��@��X�uҋT$(;�}$�D$�|$ ������ ���D����;��\��|�D$���҉T$(������T$,��;U�T$,�n����|$0�E(��t�L$<��L$8��T$$R�U������_^[��]�$ _^��[��]�$ �I �����HS�\$P3���V����   9F��   9F��   �L�W�����D$\�����$�   �D$,+ˋ�P�~8����V�T$@R�L$,�,���P�L$�2����L$������u*�D$P���	Z ��u��t��Bj����_^3�[��H� ��_^[��H� �A������������̋D$� �T$�D$V�t$ ����D$�������A��@���B�����A�^�H��B�����A�^^� ��j�h�d�    PQV�  3�P�D$d�    ��t$賶���N�D$    �T4�m����ƋL$d�    Y^�������������鋶�������������V���P4�҅�3�^�SW3��   ���������   �҅�t��u�؃�����|�_��[^�_[3�^���SV��~ Wt
�~ t��2��D$�D$ �|$$��D$��~ t�N�P���   ���$�Ѕ�u2���؃~ t$�N�D$����   W���$�Ѕ�u_^2�[� _^��[� ���������������SV��~ Wt
�~ t��2��D$�D$ �|$$��D$��~ t�N�P���   ���$�Ѕ�u2���؃~ t$�N�D$����   W���$�Ѕ�u_^2�[� _^��[� ���������������j�hX�d�    P��0SUVW�  3�P�D$Dd�    ��|$T����   ��PlW�L$Q����3�S�L$�\$P�K����5��l$X����Dz6j�L$�-����5�����Dz�E �M�U�D$�E�L$�T$�D$ �L$$������RlW�D$8P���D$T��PU�L$,�D$T腶���L$4�D$L��  �L$$�ޟ�����L$$u2�\$L�}�  �L$�D$L�����l�  3��L$Dd�    Y_^][��<� S�~���S�L$���r���� �] ����DzIj�L$(�[���j�L$���N���� �] ����Dz%�L$$�\$L��  �L$�D$L�������  �   냍N(���  ����!���L�����   �T$$R�ЍL$$���\$L��  �L$�D$L������  ���:�������j�h��d�    P��SVW�  3�P�D$ d�    ��|$0��w>����   W�҅�u/��PlW�L$Q���҃|� �D$(    u(�L$�D$(�����1�  2��L$ d�    Y_^[��� �L���T$4���   R�Њ؄�t���� ���N(��  �L$�D$(�������  �ËL$ d�    Y_^[��� ����������j�h��d�    PQ�  3�P�D$d�    jX�4�����D$���D$    t�������L$d�    Y���3��L$d�    Y���������������j�h�d�    PQVW�  3�P�D$d�    ��jX�D4�����D$���D$    t���������3����D$����tW��� ����ƋL$d�    Y_^���������������VW�|$��t5hpd���� ����t%�t$��thpd��� ����tW������_�^�_2�^�������������j�h#�d�    PQV�  3�P�D$d�    ��t$��2�D$   �u����N(�D$ �8�  ���D$������: �L$d�    Y^�����������j�hS�d�    PQV�  3�P�D$d�    ��t$�C: �N�D$    ��2�-����N(�%�  �hd���D$t��D$P���F    �F    �����ƋL$d�    Y^��� ������j�h��d�    P��   SUVW�  3�P��$�   d�    ��$�   �վ����P43ۋ�3��\$��;ǉD$�D  �L$l������L$@��$�   �����FPƄ$�   �|$�����؃�;�u0�N݄$�   ����   W���D$x�$P��;ǉD$��   �\$l�FP�   �Ӽ��������u*�N݄$�   ����   P���D$L�$P�ҋ��~�|$@��tm��ti�L$ �����D$��V�L$,Ƅ$�   �D$(蒡����$�   �L$ QWS���������u	���½����D$;ŉD$}�l$�L$ Ƅ$�   诮���L$@Ƅ$�    �.	���L$lǄ$�   �����	���D$��Ë�$�   d�    Y_^][�Đ   � ������j�h��d�    PQ�  3�P�D$d�    jX�0�����D$���D$    t�L$Q���i����L$d�    Y���3��L$d�    Y����������V��������D$t	V�[2������^� ��j�h�d�    P��SUVW�  3�P�D$$d�    ��t$4����   �E �PlV�L$Q�����D$8j��3��$�ȉ|$8�a������L$���D$,������  ����   �D$@� 3ۅ�tP�����������ty������O(��  �L$D���tP�����؃���tQ���Y���K(�q�  ��uU���������;�tU���T�����uU�z��������;�tU���7���;�u;�u>3��L$$d�    Y_^][��� �4�   �>��t	��Bj��;��>    t"�t$4�4�   ���t	��Bj���    �.�D$8����   �P�V���$�҅��D$@u9�8 u��t��Bj���ЋL$D�9 �]������U�����Bj�����E����8 u�8�D$D�8 u��   �+�����������V�t$��th`e���;�����t��^�3�^���������������̸`e�����������VW�|$W��������~ t�N��P0W�ҍNh���  _^� ����j�h9�d�    P��V�  3�P�D$$d�    ��t$�5 h(��L$�D$0    ��4�F    辝���D$Ph�=�N��  �H+���\$�N@���D$<�$�]����H+���\$�NP���D$<�$�>����Nh�D$,�F`    �z�  �Xe��t��ƋL$$d�    Y^��(������������̃�VW�������N��t��Pj���F    h(��L$������D$Ph�=�N�M& �H+���\$�~@����$衦����W�G�NP�O�VT�FX�N\_�F`    �Nh^���v�  ������VW������ ��t�O��P�����_^���������������V��~ t�N��T$�@R����D$�NQj0P�Ƅ �V@RjP躄 �NPQjP讄 ��`VjP袄 ��0^� �����������SU�l$��;�tp�����U���H �M��t�����CVW�u�{�   �E@�C@�MD�KD�UH�SH�EL�CL�MP�KP�UT�ST�EX�CX�M\�K\�U`�uh�{h�   �S`�_^]��[� �������������U������4SVW��� u �E��th7P��)����3�_^[��]� �O��u�PV�҅�u��t�h�6V�)����3�_^[��]� �O��P4�҃�t��tPh�6V�)����3�_^[��]� �O�� ��u��t�h�6V�e)����3�_^[��]� �_@���͓����u;��t,j��謒�����$j ��蝒�����$hP6V�)����3�_^[��]� ���7����T$8�H6������z0��t���$h 6V��(����3�_^[��]� ��3�_^[��]� ����������;����Az'��t�D$8���$h�5V�(����3�_^[��]� ��P���������u?���X���j���ؑ�����$j ���ɑ�����$hx5V�H(����3�_^[��]� _^�   [��]� ������������V�t$WV���������'���` th�7�h�7V��'����Sh�7V��'�����GP���*��h�MV��'�����O(Q���*��h�&V�'�����_@j���������$j ���������$ht7V�'�����_Pj���������$j ���Ր�����$hD7V�T'����� [t'h87V�?'�������&���O��BV�Ћ���&������&��_^� �������V�t$Wj ��j����*������tj�GP���[I���O@Q���`J���WPR���UJ���GhP���:I���O`Q����$��� ��t!j��"������t�WR������_��^� j �"����_^� ������̃�SV�t$W���D$P�L$3�Q�Ή\$�\$�\$�u*����;��X  �L$����   U�WR���a���o@U���v���GhP���K���O`Q���P���T$R������|$ ��t?�D$ P���D$$    �F����؋D$ ��t!P��������Gu�L$ ��t	��Bj�ЍwPj �������͋������j��������͋��b����]_^��[��� ����   �OQ������W@R������GPP������OhQ������W`R������D$P�����8\$��t=�L$Q�Ή\$ �������D$;�t!P������;ÉGu�L$;�t	��Bj�Ћ�_^[��� ��������́��   SUV���P0Wj�ҋ�$  S�������N��t��PDS�ҋ��3�L$@�.����L$(�%����L$�����D$X�~P���] ��L$�P�T$�H�L$�P�T$�H�L$ �P�D$P�L$D�T$(趑���L$@�-����L$@Q�T$R�D$`P�I�����L$4�P�T$8�H�L$<�P�T$@�H�L$D�P��S�ωT$@�U ��u3�D$pP���� �L$p芛����$����Dz�L$Q�T$\R��������D$@P��$�   Q���"���T$(R��$�   P���"����$�   Q��$�   R�D$`P蘝�����L$pQ�L$\�'�����$����zB��$�   R��� P��$�   P���˕����N(�P�V,�H�N0�P�V4�H�N8�P�V<�~h���N�  ��$�   P���oE ��   󥍌$�   ��  _^��][���   � �����������U������t  ��SV�\$|��W�L$P�t$D�D$7 �7����~` t)�E�E$���E�]�]u	�E$   ���u�E$   �^@�~PS���������t?��^X����D{3�FH���#���FX�'��ݜ$�   �E�$����������$誋���]�E�x �\$8�E�Cy �D$8�~ ݔ$�   ����ݔ$�   ����ݔ$�   ݜ$�   ��ݔ$   ݜ$�   ݜ$�   ݜ$�   ��  �N��P4�҃��D$8t	���o  �M$���3���w�$��4�   �����N�E�u(�}�]�V�u P���   VWS���$�Ѕ������D$7�  �L$D��$�   ��R� ��$�   ������L$h踑����$�   P��$�   脎����$�   �������$�   Q��$�   R��$  P�������L$t�P�T$x�H�L$|�P��$�   �H��$�   �P���|$8�ÉT$|�D$(��  ���  ���׍։T$,�P��׍։T$8�P����������ǍK��������ƉT$0�D$H�A���+������T$,������\��\$,���B�\����D$(�+T$H������ǃ�\$H�\�����B�\��A��D$(�+T$0������ǃ��l$(�\��\$0���B�Q��\��A��+T$8������ǃ����\�����BӃ|$(�\��T$8�5����D$(�]��|R������ɉL$,���ύX�ΉD$8��C�Ù+������ǃ����\�����AL$,�l$8�\�u΋]�؋D$D��P��$  RV��$,  �U�����螑��P�L$T�t�����$�   P�L$T賑����L$hQ�L$T裑���^��$�   R�L$T菑���^����   �   �\$8�A�D$H���+������ߍ�P��$$  �D$4�ϓ���L$P� �\$P�@�\$X�@��$�   P�\$d�*����L$0�T$h�R�L$T�������ލ�$�   P�L$T������\��l$8�L$H�r����]�ۋˉL$(�.  ������  ��������D$,�A���+�����ǍL��D$0    �L$8�  �����#  ���׍T��T$0�P��׍T��T$8�K�P������ۍ��������ǍT��T$,�T0�T$H�A���+����T$0�����B���\$0�\������B�\����D$(�+T$H�����B��ǃ�\$H�\������B�\��A��D$(�+T$,�����B��ǃ��l$(�\��\$,����B�Q��\��A��+T$8�����B��ǃ����\������BӃ|$(�\��T$8�)����D$(�]���s���������ɉL$,���ύX�L��D$8��$    �A��C�Ù+������ǃ����\������AL$,�l$8�\�uˋ]�����I �D$H�K�A���L$0�+������ǁ�  �yI���A;\$(݄��   ��݄��   ����܌$�   �\$H�������L���ݜ$�   �����L���ݜ$�   }����D���$�   R����$,  �$P�َ��݄$�   ��P��$  Q�T$pR����$|  �$P讎��݄$�   ��P��$\  Q��$�   R����$T  �$P耎������覍����蟍��P�L$T襌���D$P�D$8�D$0�X��D$X����D$`�XD$,�ۉD$8������L$(��؃��L$(������]�D$D��@��@�F�^�@ �F�^�x` ��   �   ;ىL$(�}   3ۅɉL$D~g�A���+����L$D��ύ���΃����D�����\�������\���D���D���\���\�������΋L$D��;��։L$D|��L$(��;M�L$(~��D$7_^[��]�$ ��}-}-�-�-��������U�������(���E��������D{�E� �$���$�H�\$��U���E��������D�E{� ���\$�@���\$�H�D$�\$ ����@�a� �a�@�E �a�A(���A �����A0�����A8���A@�������IH�����IP���IX���A`��������B���������������������A ���A�A8�����AP������A(���A�A@�����AX�����X�A0�����A���IH���I`���X���]� ���������������j�hh�d�    PQV�  3�P�D$d�    ��t$�s����N�D$    ��7�-����N �%����N8�����NP�����ƋL$d�    Y^�����V���8����D$t	V�������^� ��U����j�h��d�    P��(  SVW�  3�P��$8  d�    ��~ �D$+�~` t�E�E�E�]�]�E�]��]�E�E����E�L$4����$hhY�0* �N@�VD���ĉ�NH�P�VL�H�P�D$<P��$�   Ǆ$T      � �~Pj��Ƅ$D  �������$j ����������$�   �$Q��$`  � �ES����$X  �$Ƅ$L  ��1 ��u�D$+�~ t$�v�E�E����   P�����$�҅�u�D$+��$L  Ƅ$@  � ��$�   Ƅ$@   �s �L$,Ǆ$@  �����?  �D$+��$8  d�    Y_^[��]� ���U����j�h�d�    P��(  SVW�  3�P��$8  d�    ��~ �D$+�~` t�E�E�E�]�]�E�]��]�E�E����E�L$4����$hhY�( �N@�VD���ĉ�NH�P�VL�H�P�D$<P��$�   Ǆ$T      �h �~Pj��Ƅ$D  �T�����$j ���E������$�   �$Q��$`  ��� �ES����$X  �$Ƅ$L  �m1 ��u�D$+�~ t$�v�E�E����   P�����$�҅�u�D$+��$L  Ƅ$@  ��  ��$�   Ƅ$@   �� �L$,Ǆ$@  ����� �D$+��$8  d�    Y_^[��]� ���U����j�h_�d�    P���  SVW�  3�P��$�  d�    ��E���.  3�9^�#  3�9^`t	�   +ȋ�;��s  �L$t�� �E�N���T$T�$R��$  �'���D$LP��$   �~Q���@ ��T$t�H�L$x�P�T$|�H��$�   �P��$�   ��$�   �@Q�ω�$�   �	 ���$�   �H��$�   �P��$�   �H��$�   �P��$�   �@�L$tQ��$   R�L$T��$�   �n������$�   �P��$�   �H��$�   �P��$�   �H��$�   �P��$�   ��$�   �G���ݜ$�   ��$�   �t������  �N��@h�T$dR����$�����$Ƅ$  ��|������$  �$Q�N������T$L�H�L$P�P�T$T�H�L$X�P�T$\�@�L$d�D$`��$   �3�  �L$LQ��$   R���	 ��$�   P��$  Q�L$T�f������$�   �H��$�   �P��$�   �H��$�   �P��$�   �@��$�   ��$�   ������u��$�   Q��$�   ������$�   R��$�   P��$  Q�z������$�   �H��$�   �P��$�   �H��$�   �P��$�   �@����$�   ��$�   � ����L$t�U���N@�VD���ĉ�NH�P�VL�H�P��$�   P��$@  �G h�   Ƅ$  ��������|$d;�Ƅ$   t1��Pj���{�����$S���{������$<  �$Q���� �3���$,  ����$   �� �L$tǄ$   ������ �ǋ�$�  d�    Y_^[��]� ��uy�N��Bd�Ћ�;�ti�E�^@�NP�\$dS袐����t"�E���NP�$�z�������$�pz���\$d���\$d����D{#�NQ��$  R� �D$hP�����$��1 �ǋ�$�  d�    Y_^[��]� 3���$�  d�    Y_^[��]� ��������U����j�h��d�    P���   SVW�  3�P��$�   d�    ���|$0�u���D$(    t	����  �]���z������  �` t	�   +Ƌ�����  �L$D�Ny����$   �wPVS�L$L������L$D�`z�����I  ���Qz�����:  ��@���?z�����(  j �L$H�y��� �����$�]y���\$\j�L$H��x��� �����$�?y���\$T�L$4��x��j �L$8Ƅ$  �x���D$\�����$�D$4��x���L$,�j�L$8�x���D$T�����$�D$4�x���T$,�L$4��Ey������;������zH�H6����Az=�D$4�L$8�T$<��D$@�O�W�G���S�V�C�F�K�N�D$(   ��؍L$4Ƅ$    ���  �L$DǄ$   �������  �|$0�Q�L$DǄ$   ������  3���$�   d�    Y_^[��]� ����   �O����   ����   S�ЉD$(�|$( tw�_h�   ��|$d��Ǆ$      �U�  ��$�   Q�L$4�t0 ��$�   �(�  ��������t�L$d�Ԋ����t�T$dR����  �L$dǄ$   �������  �D$(��$�   d�    Y_^[��]� ����U����j�h�d�    P���   SVW�  3�P��$�   d�    �ً}��t	���(  ����   W�҅��  �D$/��PlW�L$8Q����j �L$8Ǆ$      �v���uj �ΉD$4�v���D$0�����z#j �L$8�Xv��j �ΉD$4�[v���L$0��D$/j�L$8�5v��j�ΉD$4�8v���T$0�����A�d  j�L$8�v��j�ΉD$4�v���D$0��{` t	�   +ϋ����D$/ �c  W�L$8��u��� �sP�����$�!v���\$\j�L$8�u��� �����$�v���\$T�L$D�u��j �L$HƄ$  �{@�u���D$\�����$�D$8�u���T$0j��L$H�Zu���D$T�����$�D$8�eu���D$0�L$D��v���H6����Au(j �L$H�u��� �H+j�L$H�\$X�u���D$T��L$D�T$H�D$L��L$P�W�T$4�G�D$8��T$@�O�L$<�F�N�L$D�V�D$/Ƅ$    ��  �\�|$/ ������L$4Ǆ$   �����d�  2���$�   d�    Y_^[��]� ��up�K��ti����   �T$4R�Є��D$/tR�������Ch�   ����$�   ��Ƅ$   ��  �L$dQ���2- �L$d���  ��$�   Ƅ$    ���  �L$4Ǆ$   �������  �D$/��$�   d�    Y_^[��]� �����3�9A`���A`�   ���������������̃y �tW�y` t�D$��D$�D$<�T$�I����   ��(�\$ �D$\�\$�D$T�\$�D$L�\$�D$D�$R�T$0���$R���@ �������������̃�V��3�9F`t3�9D$����L$��uZW�N�G� �~@j ���s��� j�\$����r��� �H+���D$�����\$���$軄���NP�v��_�   ^��� ��u9Ft�N����   ��^��� ��������U����j�h1�d�    P��(  SVW�  3�P��$8  d�    ��}3�9F`��;��2  ����$�L$4hhY�C �N@�VD���ĉ�NH�P�VL�H�P�D$<P��$�   Ǆ$T      � ��Pj��Ƅ$D  �r�����$j ����q������$�   �$Q��$`  �� �E$��Ƅ$@  t���3��E4�U(�M���\$�E,�$R�EP�E P���\$�E�$Q��$|  �o����$L  ��Ƅ$@  �� ��$�   Ƅ$@   � �L$,Ǆ$@  �����Q �Ë�$8  d�    Y_^[��]�4 �E$��t���3��E4�N�u(����   ���\$�E,�$V�EP�E P�E���\$�E�$P�ҋ�$8  d�    Y_^[��]�4 ������̃�`SV��L$2���w���L$ ��w���D$l����   �~` t��w�$��H����   ����   �L$PQ�N�����T$�H�L$�P�T$�H�L$�P�T$�@�L$Q�T$TR�N�D$$�� ��L$ �P�T$$�H�L$(�P�T$,�H�L$0�P�D$ P�L$Qj j�T$D聛 ����^��[��`� �N�D$8P����g���^3�[��`� ��H�G�H�H����V3�9q`t3�9D$����D$��u��@�]p����7����u$�   ^� ��u9qt�I����   ��^� ��^� ������j�hk�d�    P��   SVW�  3�P��$�   d�    ���P3�W�҅�t�D$(P�N�� P�L$Q�N���P�L$H��M��݄$�   �N����   ���D$H�$P��$�   �ҋ؅�t��$�   ��t�    �t$@�L$@Ǆ$�   �����i�  ����ǋ�$�   d�    Y_^[�ļ   � ��������V3�9q`t3�9D$����D$��u��@�o����7����u$�   ^� ��u9qt�I����   ��^� ��^� ������W3�9y`t3�9D$����D$��uNV�qP���
o����tt�D$�D$�L$PQ���$j����m�����$j ����m�����$�o� �� ^_� ��u*9yt%�D$�D$�I����   P�D$P���$��_� ��_� ^��_� �����������SV��2ۃ~` t�   +D$��D$��u:�D$�D$������zh�����\$�NP�$��~����P0j���ҳ^��[� ��u>�~ t8�N�D$��Pl���\$�D$ �$�҅���P0j������^��[� ����^��[� ������������j�h��d�    P��VW�  3�P�D$ d�    ���D$    �t$0���D$(    �^l���` �D$(    �D$   t�   +D$4��D$4��u�GP��OT�N�WX�V�G\�F�9��u4� t.�O��Rh�D$P�ҋ��P�V�H�N�P�L$�V�ú  �ƋL$ d�    Y_^�� � �������������U����j�hءd�    P��   SVW�  3�P��$�   d�    ��3�9F`t�M�]���}��]�}9F��  �N��@h�T$DR�Ћ�����3���$�   �D$0����L$l����T$p����D$t����L$x�L$T�T$|��$�   �Gr������T$<u���  3��\$4�|$,�D$,�L$0Qj ����T$\R���L$X�$��j���N���$��������   �L$T�T$X���ĉ�L$t�P�T$x�H�L$|�P��$�   �H�N�P�7� �D$4������z�\$4���h���L$p��s����t�D$TP�L$p�����D$<�\$<�L$T�T$X�D$\�L$l�L$`�T$p�T$d�D$t�D$h�L$x�T$|��$�   ����@�|$,������t�N@��j���L$4��E��t
�D$<���؍L$DǄ$�   ����蠸  �   ��$�   d�    Y_^[��]� ����t���t���$�   d�    Y_^[��]� �؋�$�   d�    Y_^[��]� ���VW��3�9~`t�   +D$��D$��uR�NP�jj����t_�N@�j�����8������u_�ظ   ^� � 8����Az
_�   ^� _�   ^� ��u9~t�N��Px��_^� ��_^� U������4SVW��3�9~`t
�   +E��E����   �^P����i������   �3�9~`����P�Bt�Ћ����|$4��   �D$4j ������\$<�h���M�   �;��t$4~&�D$4�����L$@�$�hh���U���;��t$4|�j���>h���E���   _^[��]� ��u9~t�N��E�R|P��_^[��]� ��_^[��]� _^3�[��]� ���3�9A`t�   +T$��T$��u�B� ��u9At�I����   ��� �����̃�h�x�  ��������j�h�d�    PQ�  3�P�D$d�    h�   �U������D$���D$    t���K����L$d�    Y���3��L$d�    Y������������j�h;�d�    PQVW�  3�P�D$d�    ��h�   ��������D$���D$    t����������3����D$����tW�������ƋL$d�    Y_^������������VW�|$��t5h`e���j�����t%�t$��th`e���R�����tW���f���_�^�_2�^�������������j�h��d�    PQV�  3�P�D$d�    ��t$��4�D$   ������Nh�D$�ش  �NP�D$�˴  �N@�D$辴  �N�D$ 豴  ���D$�����B �L$d�    Y^����U����j�hܢd�    P��h  SVW�  3�P��$x  d�    �ى\$43�9{�|$8��  ��$P  ������$  ��$�  �ڦ����$�  Ƅ$�  �F� h(�h�=��$�  Ƅ$�  �H@����s@ݜ$,  j���#e���\$<W���e���l$<����$�  �$�1� ��$P  P��$�  ��	 ���  �{P����e����t*j����d�����$j ���d������$`  �$�����K�E����   j ����$  �$P�҅��D$8��  ��$  u*hl8hP8hd  h48�X����j��$  轢����$  tuh8hP8hi  h48�W������$�  Ƅ$�  �3� ��$  Ƅ$�   �������$P  Ǆ$�  ���������3���$x  d�    Y_^[��]� j ����c����$����D{-�KQ��$8  P��� Pj ���c������$  �$�+ ��$�   �/����K�S�C�{��$�   �O��$�   ��$4  ��$�   �W��$�   �GQ��Ƅ$�  ��$�   ��$�   �y� ���$�   �H��$�   �P��$�   �H��$�   �P��$�   �@��$�   ��$   �bq����$�   Q��$�   ��f����$�   �Bq����$�   R��$�   P��$<  Q�Us�����$�   �H��$�   �P��$�   �H��$�   �P��$�   �@����$�   ��$�   ��p���u��$�   Q��$  R��$X  P��虠����u��$�   Ƅ$�  �w���������$|  Q��$  ������$�  R��$  �$�����$�   �i���L$l��h���L$L��h���5�D$D�T$DP�\$@��$�  Q���4� ����   �D$D���$�Ma��������   �D$D����$<  �$R���	� � ݜ$�   ��$|  �@ݜ$�   �@��$�   Pݜ$�   ������;����AzY3�9^~N�d$ j S���fW���T$d݄$�   �L$L��Qj S�\$X��݄$�   ���\$`܌$�   �\$h��q����;^|��\$4�T$<R��$�  P���N� ����   �D$<���$�g`��������   �D$<����$<  �$Q���#� � �\$l�T$l�@R�\$x��$�  �@ݜ$�   �����;����AzW�^3���9~~F�SW���V���T$d�D$l�D$L��PSW�\$X��݄$�   ���\$`܌$�   �\$h�q����;~|��\$4�{` t����   ���Ѝ�$�   Ƅ$�  �Au����$�  Ƅ$�  ��� ��$  Ƅ$�   ������$P  Ǆ$�  ��������3�9D$8��������$x  d�    Y_^[��]� �����������U����j�hS�d�    P��(  SVW�  3�P��$8  d�    �L$D�E�3�;މt$`th`e���������u3ۋM�9;�th`e���������t�|$H��t$H��;�t;�u3���$8  d�    Y_^[��]� �U92t;�tۋE90t;�tЋE;�t��uċ|$D9w`t
�   +ȉM�L$t�t$L�t$P�l^���L$d��$@  �\^����$�   Ƅ$@  �H^����$�   Ƅ$@  �4^���GD�W@�OH�t$D��@�D$x��T$t�W��P�D$d�G�L$|�O��$�   �W�D$p�F�L$h��T$l�V��$�   �F��$�   �N��$�   ���$�   �E����$�   �N��$�   �VƄ$@  ��$�   ��$�   �  �E�����$��]���\$T�Ej�����$��_������  �D$T��$����A��  ��������A��  �����$�`]���T$Tj�����$�_�����}  j�L$x�D$d   �]���D$Tj ��L$h�]���D$Tj���$�   ��\���Ej ���$�   ��\���E�t$D�;�u�F��N����9t$H�N�D$Lu	�L$P�   �����D$P�   ����  �t$D�~ ��  �N�E����   �D$PP�D$PP���$�҅��D$`��  ;�u�N��t	��Pj�ҋD$L�C�!�|$H;�u�΋I��t	��Bj�ЋL$P�O��h�   ��$�   ��Ƅ$@  uPh�   ��������D$T��Ƅ$@  t��������U�|$DƄ$@  �؉�6�U�|$D3�Ƅ$@  �؉��|$D;�t�K��t��Pj���C    �t$H��u;h�   �m������D$T��Ƅ$@  t	���c����3��MƄ$@  �D$H���;�t�N��t��Bj���F    �w�{�   �L$t�K@�T$x�t$D�SD�D$|�CH��$�   �KL��$�   �SP��$�   �CT��$�   �KX��$�   �S\�F`�C`�L$L�K�Kh�L$T蠩  �D$H�x���   �T$d�P@�L$h�HD�T$l�PH�L$p�HL��$�   �PP��$�   �HT��$�   �PX��$�   �T$D�H\�J`�H`�T$P�ph�ΉP�0�  ��$�   P���Q ��$�   ��  �|$T���m����t��$�   �m����t��$�   Q���W�  �L$H��$�   R� ��$�   躨  ���sm����t��$�   �cm����t��$�   P����  ��$�   Ƅ$@  �|�  ��؍�$�   Ƅ$@  �d�  ��$�   Ƅ$@  �P�  �L$dƄ$@   �?�  �L$tǄ$@  �����+�  �D$`��$8  d�    Y_^[��]� ���������������V��������D$t	V��������^� ��U����j�h��d�    P���  SVW�  3�P��$�  d�    ���|$�Oh�`l���Ѕ��  ��$4  ��  ��$d  Ǆ$       �Ҧ  ��$  Ƅ$   辦  �Oj ��$h  PƄ$  � ���D$�c  �L$�_����L$Q��$h  Ƅ$  ��  �L$,�m_���L$D�4� ��$�   �ORƄ$  �� ���$�   �P��$�   �H��$�   �P��$�   �H��$�   �P�w@j�Ή�$�   ��W��ݜ$�   j ����W��ܬ$�   ���L$L�$��� 3ۋD$ ��L$,�T�T$0�L�L$4�T�T$8�L�L$<�Tj �D$0P��$  �T$H��  ��$�   Q�T$0�wR����� ����  j�D$HP��$  ��  ݄$�   ����$�   �$Q���� ��T$D�H�L$H�P�T$L�H�L$P�P�T$T�@�L$DQ��$�   R�L$4�D$`�
`����L$\�P�T$`�H�L$d�P�T$h�H�L$l�P�L$\�T$p��d��ݜ$�   �L$\�(e������   ��$�   P�L$`��_�����5����A��   �L$\Q��$�   R��$�   P�g�����$�   �P��$�   �H��$�   �P��$�   �H��$�   �P���L$t��$�   �d����th�L$D�N0����$�   Pj �O@��U�����L$P�$�:���L$D�t� ��t1��$�  Q�L$H��� ��   ��$  󥍌$�  �s�  �|$��$  R��$8  諧  �����   �������$4  � i����t��h�   ��$4  �|$�D$   �L$DƄ$   �n� �|$( Ƅ$   �D$�$t"�D$ ��t3�VP�L$$��$�t$ �t$(�t$$��$  Ƅ$   ���  ��$d  Ƅ$    譣  ��$4  Ǆ$   ����薣  �|$ ��   �T$�M�ɋutH��t3��_h����Au�Gh��A�_p����Au�Gp�Y�A�_x����Au��Gh��Gp�Y�Gx�Y�M����   ��tc�ܟ�   ����z݇�   ��Aܟ�   ����z	݇�   �Y�Aܟ�   ������zY݇�   �Y��$�  d�    Y_^[��]� ݇�   �݇�   �Y݇�   �Y��$�  d�    Y_^[��]� �D$��$�  d�    Y_^[��]� ���V�t$��thPf���k�����t��^�3�^���������������̸Pf�����������U����j�h�d�    P���   VW�  3�P��$�   d�    ��$�   �SZ���L$d�JZ���L$L�AZ���L$|�8Z����Ph�L$<Q����j �L$@Ǆ$      ��R��� j j ��$�   Q��$�   R�����$��������  �L$|�@a�����  �D$|P��$�   Q��$�   �[����T$d�H�L$h�P�T$l�H�L$p�P�T$t�@�   �D$x�t$4�   ;��|$0��   �D$4�\$4�D$0���L$D�t$<�$�MR������$�   �$Q���X�����T$L�H�L$P�P�T$T�H�L$X�P�T$\�@��$�   Q��$�   R�L$T�D$h�[��P��$�   P��$�   Q�M��0����uJ��;��|$0�f��������t$4�=����L$<Ǆ$   �����V�  2���$�   d�    Y_^��]ÍL$<Ǆ$   �����+�  ���$�   d�    Y_^��]�����U�������   ����� ���@  ���� ���1  ���/� �\$H���$� �T$P�D$H������u�������������u���T$8��T$8������������  ��������  ��'������A��  ����'�T$p������������A��  �������������]����A��  �D$XP����� P��$�   Q���� ���	o����;�������O  �D$8�p&�������:  �WHR�NH�sY���\$8��8�< �T$@�D$8��������t�E������A{�xD����{2���]��؋���V��P��$�   P��$�   Q���q� ����X������V��P�T$|R��$�   P���� ���X����$�   �^���L$x�^���L$xQ��$�   ��X���D$@������A{�E������A{�xD����{2���]��؋��� ����\$@�� ���T$8��$�D$@������Au�����T$@��������Au���T$8������D$H���D$P����������Au�������T$@���������z�������\$8�������;����������   ����������A��   �N< �L$H�\$X�D$8�=< �L$P���l$`�$�D$H��: ���d$P���\$`�D$@��: �D$X�%�$���L$h���D$h�$�c���L$X�X����;������z#�\$p����Au���]�����2��؋�]���������2���]����������������U����j�h1�d�    P��  SVW�  3�P��$�  d�    ����~ �  �V���  �^;���  ��|D�F�L���A�Y����Dze�A�����DzL��Y�����DzE�A��Y�����Dz=���� ��Å�~1�N����    ��Y�����Dz�����������������J�;��p  �C�;��e  �F���������Q  �F�D��������A�<  �F��D��������D�%  �F�N��+؃���D��������D�  �F�V�L8���D��������D��  W���>p����$����D��  �L$(�č���F�N�V�D$8�D$<�F �D$H�ÉL$0�T$4�V��    ыN(�T$D���L$TǄ$�      �T$P��� ��;���L$0�$Ƅ$�  膓�����   ��;���$�D$\Pj �L$8�Rz������   ��$�   �� ��;�V �N�׍�    ȋF(�L$D�ЉL$P���L$0Ƅ$�  �$��������   ��;���$��$�   R�D$`P�L$8��y����tq�E���\$��$�   �E�t$d�$���������tJ��Ƅ$�  �-� ��Ƅ$�   �� �L$(Ǆ$�  �����ں�����$�  d�    Y_^[��]Í�$�   Ƅ$�  ��� 3��L$T�D$D�D$P��$�  ��� �L$(Ǆ$�  ����耺��2���$�  d�    Y_^[��]���������U������t  SVW��3ۍ�$0  ��$�   ��$�   �cQ����$H  �WQ����$�   �KQ����$�   �?Q����$   �3Q����$  �'Q����$�   �Q����$�   �Q���L$h�Q���L$P��P���u ;�u
��$�   �u �U$;�u
��$�   �U$�E;�u
��$`  �E�M��u2�_^[��]�0 ��u4�E0���\$�E(�$R�EVP���\$�E�$Q���G���_^[��]�0 �E�]����D{��Q�5�������Q�L$P�����؃����]t
��t��u�~���D$?t�D$C��D$? ���D$C �D$B u�D$B�O3�8D$?�D$H   ����+����D$Du�D$D    �E�E��������Au�����   �R�WP�G���$PRQ�2� �O���D����������������@� ������4u��D$@}�D$@ �E�_�E�D$A �эT3�������  �T�����zV�D���������zM�D�����������Az>�O�B;�}4�G���D��U ��URj���$PQS�~� �E�����������ـ|$@ ��&t�����T$���$V������E�D$A��؋E �0�O�_�t��K���+փ�|;�G�T��R�����uV�R�����u?�����u;�R����u6���A��� ;�|�;�}0�W�������u����;�|����������;���  �T$L;Ut[�G�T���L������zI��E��������u7�E0�M$�E ���\$�E(�$Q�MPQ���\$���$R����_^[��]�0 ��2���_^[��]�0 ������AuR����������AuJ���$���������Az<�C�;�~5�����ЋM ��URj����$P�GPS�� �E�����������ـ|$@ ��&t�����T$���$V�@����E�D$A��؋] �3�G�t��H���+у�|;�G�T���R����AzV�R����Az?�����Az;�R�����Az6���A�� ;��;�~,�W�������Az����;�����������;�S�T$L;U������G�ȍ�����A�������E��������������E0�M$�E���\$�E(�$QSP�p����L$D���D$H�����L$D�E������u��ݔ$�   ��ݜ$�   �ݔ$�   ��ݔ$�   �ɋ_��������   ݄$�   ������A��   �|$H ��   �G�P���+ƃ�|F�O�L��A��Y�����Dza��Y�����DzH�A�����DzA�A�Y����Dz9���B��� ;�|�;�}3�O���A�����Dz����;�|����������;���   �L$L2�;M�����E0�E$�U ���\$�E(�$P�E�ERP���\$�$Q�������_^[��]�0 �G�P���+�|F�O�L���A�Y����Dze��Y����DzL�A������DzE�A��Y�����Dz=���B�� ;��;��Z����O���A������Dz����;�����������;��'����G�T$D���������D��  �}���  �|$? ��U Rj�tX��$  P��$�   Q��$@  R�����$������E Pj��$   Q�O��$�   R��$X  P�����$������F��$�   P��$<  Q�����$������U R�W��j��$�   P��$T  Q�����$�����|$B �u  �\$C��tL�D$hP��$�   Q��$  R��$�   P��] �L$`Q��$�   R��$0  P��$�   Q�] �� ��   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��O����$�   ��O����$�   R��$�   �J���E(��������A�	  ����  �E0�L$P�T$T�]��(�\$ �ă����\$0���$�   �P��$�   �H��$�   �P��$�   �H��$�   �P��$�   �ĉ��$�   �P��$�   �H��$�   �P��$�   �H�Pu�A�����*�����@���  ��u$�E0���\$���E(���$����������   �|$@ �  ��&���|$X �T$�$}��+G��P�	��+O��Q���Y���8D$A��   �E$�U�    �O���_^[��]�0 ��$�   �DM����4����$�   �$R��$t  P��$�   ��H�����O������   �|$? t`��$   ��L����4����$   �$Q��$t  R��$  �H�����;O����u!�E$�U�    �O���_^[��]�0 ���Et$H�_��ܜ$�   ����A�	����X����؋E$�U�    �O��_^��[��]�0 �U������4SV��~W�D$;�EP�����������U�F�N�D���E��������A��  �F�T��������  R���.����N�V��;ʉE�l  ���c  �} u�D$<�D$<    �E�E�E� P�Fj���$PRQ�� �^�ЋF�L��D��<������������@� �F��������4� ���@��������Auc�E���'��������Az�C�;�~������]�A�g��������Az3�~�A;�})�F�D��M��URj���$PWS�l� ������؅�}3ҋE��F�|����;��h  �V�J�;��Z  �N�E������D�F  �}u2�_^[��]�8 WQR�VR�׊ �M�؍A�����
w8���|�$��|�V+Ӄ�| �_^[��]�8 �F+Ã�|�_^[��]�8 �E8�U��(�\$ �E0�\$�E(�\$�E �\$�E�$R�E���$Q���������D$;��   �}��   �F�H�;���   �P�;�~|�N��;�}r��&�����T$+��$��R��������&�؋F����T$���$+ȃ�Q������:�u$��u%�E8���\$���E0���$�j�������t�D$; �D$;_^[��]�8 �E8�E��(�\$ ���E0�\$�E(�\$�E �\$�E�$P���$R�����_^[��]�8 �L{7{a{  ��������̋L$�ɋT$�tV�D$������zG�D$������Au8������� {}������������u�����������������u	���������2�����������4�T$���$�A�D$P�D$RP���$�g���� ���̋A��3҅�~#SVW��q���<����q�<�����;�|�_^[�SU�l$VWU��萁���^3���~$��$    �F����t;�t��B0U�Ѓ�;�|�_^][� ������������SUVW��襽���N$�V�^�� �J3��ۍ,�~�V����t	��P����;�|�_^��][������������̋D$SVW���_3���~�O����t�P�B�Ѓ�;�|�W �O��Q�RP�* ��_^[� �������̋D$S��;���   UVWP�����k�{3���~����t��Pj����    ��;�|�|$�CP�O�����{$ �s|�F    �O Q���s!���F��t�N��~��    Rj P� ����P��W����_^]��[� ������������U����j�hp�d�    P��hSVW�  3�P�D$xd�    ����Ph�L$4Q�����E���\$3��E�L$4�$��$�   ��M���L$$Ƅ$�   �:����;�t$ ty�D$$P�L$8��N����tg�G ;ÉD$~Q���$    �G��    �����L$<�$��8���w��    ���L$,�$��8�����;\$|��t$ ��B0j���ЍL$$Ƅ$�    ��  �L$4Ǆ$�   ������  �ƋL$xd�    Y_^[��]� �SUV��W�}����3���~#�E����t��D$�RtP�҄�u2ۃ�;�|�_^]��[� 2҃yu3�A�8 t+��D$�T$����   ���$R�T$R�Ѕ������ ��� ��������������̋D$��@���%  �Q��;��  �I��V�0��W�x��   ����   �T$0R�������D$P��������L$Q�T$4Rj j�b ������   V�*� W���"� ������u����   ����;�\$t�N��� ܎�   � {�����T$t1�O���� ܏�   � {�D$������;����Au
�\$��������T$����Au�\$��؍D$P�L$4�;U���\$����Au
_�^��@� _2�^��@� 2���@� ���̋D$��SVW��| �{�p;�}�F�P��������u��;�|�_^3�[� _��^[� ��̋D$��|;A}	�I��� 3�� �����QV�t$W�����D$    ��5���D$��|;G}�O����W�D��^_��^Y� �VW��3�9~~C�F���t:�|$����ĉ8�|$(�x�|$,�x�|$0�x�|$4�x�|$8�x���   �Ћ���������_^� ����V��NW�A�3���|H;�}D�N����t:�|$����ĉ8�|$(�x�|$,�x�|$0�x�|$4�x�|$8�x���   �Ћ���豸����_^� ����������U����j�h��d�    P��   SVW�  3�P��$�   d�    ���|$8��Ph�L$DQ����3��L$D��$�   �5������   �_�}���t$<t\���5������   V���[I�����L$P�$�6������   V���I�����L$P�$�6������   ��T$D�G�T$L��D$D�D$L��|J�D$8�P�J������Q�������   �����uy�Q����ut�Q����uo���C��� ;�|����;�}�L$8�Q�L������uI����;�|����؍L$DǄ$�   �����S�  3���$�   d�    Y_^[��]� ��������;���}��L�������Az����;�|��;��؉\$@}��L$X�t��Ƅ$�   �ދT$8�E�B�<� ���  j ��;��$uB���}���   W�Ѓ��D$<�	  �L$8�Q�D��ڋ���\$��� �Bl�$���i� ����   �L$dQ���ҋ�����   9|$<}�|$<�D$8�H�D��ك��\$�L$h� �$��^���M�T$XR�ӧ�����L$X��   �ru����;\$@�%����L$XƄ$�    �4����E��t�M�P���   �ЍL$DǄ$�   �����ۀ  �D$<��$�   d�    Y_^[��]� �L$X��Ƅ$�    �ܡ���@����L$XƄ$�    �ơ��륍L$XƄ$�    賡���L$DǄ$�   �����o�  �ǋ�$�   d�    Y_^[��]� Ƅ$�    �x�����������SW���_��u_3�[�UV3��۽   ~2�I ��|2;w}-�G����t#����   �Ѕ�t��u���;�|�^��]_[�^]_3�[����U����j�h�d�    P��hSVW�  3�P�D$xd�    ��F �E�N�~���$PQ3���M ����}3��;�|�G����  ;F�  �N�<����  �V�D����\$�L$D� �$�WE����Ph�L$$Q��Ǆ$�       �ҍD$$P�L$8Ƅ$�   �xF���E��t^���L$<�$�0�����L$,�$�C0���]����   S�����$�Ћ���t<����L$,�$�V0�����L$<�$�0�����E����   P�����$�ҋ��L$$Ƅ$�    �~  �L$4Ǆ$�   �����v~  �ƋL$xd�    Y_^[��]� �ËL$xd�    Y_^[��]� ��������U����j�h�d�    P��hSVW�  3�P�D$xd�    ��F �E�N�~���$PQ3��'L ����}3��;�|�G����  ;F�  �N�<����  �V�D����\$�L$D� �$�C����Ph�L$$Q��Ǆ$�       �ҍD$$P�L$8Ƅ$�   ��D���E��t^���L$<�$��.�����L$,�$�.���]����   S�����$�Ћ���t<����L$,�$�.�����L$<�$�g.�����E����   P�����$�ҋ��L$$Ƅ$�    ��|  �L$4Ǆ$�   ������|  �ƋL$xd�    Y_^[��]� �ËL$xd�    Y_^[��]� �������̋T$3���|;Q}�A����    � U����j�h��d�    P��   SVW�  3�P��$�   d�    �����   �҅��]  �F���Q  ��Ph�L$dQ���D$ ��j ��Ǆ$�       �7-���Mj ���;-�������z��2ۍL$dǄ$�   ������{  ����  �~ ��  �F�8����  j �L$HQ���������Rh�D$$P��Ǆ$�      �ҍD$$P�L$HƄ$�   �<C�����Mj t�,���#�,�����L$L�$��,�����L$,�$�,��j�\$�L$(�j,��� ���\$�L$t�D$$�$�1A������   �D$dP��Ƅ$�   �҄��D$��   ��Ph�L$tQ���ҍL$dQ��Ƅ$�   �B���L$t��Ƅ$�   ��z  ��t�M�~j ��+����U��Rh�D$tP���ҋ~j ��Ƅ$�   ��+��� ���L$,�$�,�����L$L�$��+����L$tƄ$�   �]z  �L$dƄ$�   �Lz  �L$$Ƅ$�   �;z  �L$DǄ$�   �����'z  ��Ph�L$dQ����j��Ǆ$�      �5+���Mj���9+�������Au��2ۍL$dǄ$�   ������y  ����  �N�A�����  ;���  �V�<�����  ���Q�D$XP���������Rh�D$4P��Ǆ$�      �ҍD$4P�L$XƄ$�   �+A�����Mjt�*���#�*�����L$\�$��*�����L$<�$�*��j �\$�L$8�Y*���D$���\$��$�   � �$�?������   �D$tP��Ƅ$�   	�҄���   ��Ph�L$dQ���ҍL$tQ��Ƅ$�   
�@���L$d��Ƅ$�   	�x  ��t�F�V�Mj�<���)����[��Ph�L$Q���ҋN�V�<�j��Ƅ$�   �)��� ���L$<�$��)�����L$\�$�)����L$Ƅ$�   	�Ax  �D$�L$tƄ$�   �+x  �L$4Ƅ$�   �x  �L$TǄ$�   �����x  �\$��t�������Ë�$�   d�    Y_^[��]� 2���$�   d�    Y_^[��]� ���SVW���_3���~!���G����thPf謍����u��;�|�_^2�[�_^�[������VW�|$��t5hPf���z�����t%�t$��thPf���b�����tW���v���_�^�_2�^�������������j�hȥd�    PQVW�  3�P�D$d�    ��t$����3�W�N�|$��8�-����F%�~�~ �~$�ƋL$d�    Y_^������������j�h�d�    PQSUVW�  3�P�D$d�    ��t$耪���\$(�~3�S�ωl$$��8�����N�C;��D$ �%�i�i�i~P�a���G;�t�;�~��    QUP�� ���ƋL$d�    Y_^][��� ���������V��N��������~ t(�F��t!�j P�B�����F    �F    �F    ^���j�h>�d�    PQSUVW�  3�P�D$d�    ���|$��8�o���D$    �]����w3�9^t�F;�t�SP�B���Љ^�^�^9^�D$ �%t�F;�tSP���%�^�^�^�͈\$ �������D$ �����T����L$d�    Y_^][��Ãy ~�A���t��B4��3���������SV��W�{3�����3���~/�T$U�l$����t�C����@8R�T$UR�к   �;�|�]_^[� ������SU�l$VWU���P�����P0j���ҋ_3�����3���~��I ��t�G����BDU�Ѓ�;�|�_^][� SUVW���o3���~�G����t��BH�Є�t��;�|�_^]��[�_^]2�[������U������0SUVW��M�3��ɈD$:�D$; �L$<~z�E�4���tP��BH���Є�uC��BL���D$;�Є�u1��j ���$j ��轳���؅�t��Bj���ЋM����D$: ��;|$<|��|$; t�U �B0j���ЊD$:_^][��]��������SUV��W�}3ۅ���3���~$��t �E���D$��RPP�D$P�҃�;���|܋�����_^]��[� ������U������tSVW����_�P4�\$0�ҋ��L$P�t$4�E+���L$8�<+������  ����  �G �K;�t�M����  PSh;Q�}  3�����   �W�<� ����   � ��]�ȋBS�Ѕ���   �O����B4�ЋL$4;���   �O�D��������A��   �|$0~�} u�W������   �҅���   ��;t$0�w����} u+�_�   ;�~��I �F�P����������   ��;�|�_^[��]� �E����  Vh�:P蔹�������_^[��]� ����  Vh�:S�o������g��_^[��]� ���a  QPVh�:S�H������@��_^[��]� ���:  ���D����$��� �NQ���$Vh\:S������ � ��_^[��]� ����   �T$0RVh,:S��   ��� ����O��    �D���T$hR�\������L$P�P�T$T�H�L$X�P�T$\�H�L$`�P�D$h�T$d��P衸����L$8�P�T$<�H�L$@�P�T$D�H�L$H�P�D$8P�L$T�T$P�j@���E��t'���$V���Vh�9P�-������%��_^[��]� �����_^[��]� �E��tVSh�9P�����������_^[��]� �������U������t���SV�5��W�=���ًC����|$D�=��P�t$D�t$\�u�L$<�T$@�|$L�=���L$T����T$X���h�;V�D$0�|$X�L$h�T$l�|$p�\��������Ҷ��3�9|$$�  �K��    �D$(��8 t3��T$hR�E�����L$8�P�T$<�H�L$@�P�T$D�H�L$H�P�6����������D$8����L$<����T$@����D$D�L$H�L$8�T$L�1����t�L$P�1����t�D$PP�L$<�>����5�K�\$0�D������\$�O� �L$<�$Qh�;V�g�������~_�D$0���$�q������t�D$0���$h�;V�5������/�L$8�0����uh�;��L$P�s0����uh|;V������h�&V����������l����S�|$(�<: �:uJhh;V�ѵ������������D$X����L$\����T$`������D$\�L$`�T$d�D���PV�ҋC�L$h�Q�������T$P�H�L$T�P�T$X�H�L$\�P�T$`�@�D$d�������|$,;|$$�����������_^[��]� ���������j�hh�d�    P��4SUVW�  3�P�D$Hd�    ���|$�\$Xj j������������   �oU����������tUj �������j ��������L$�<l  �D$P���D$T    �����L$���D$P�����l  ��t��W���U�����3���~-��t)��|�D$;x}�H���3�P���9~����;���|ӋƋL$Hd�    Y_^][��@� �������j�h��d�    PQVW�  3�P�D$d�    ���D$    �|$ ���D$    �0���N���D$    �D$   ~2�F �Q;�u(�F�������Au�v�΃��\$����$��.���ǋL$d�    Y_^��� �SUV��W�{3�3���~"�C�<� ��t���Bx�Ѕ�t���;�|�_^��][�_^]3�[����������������U����j�h�d�    P��hSVW�  3�P�D$xd�    �ى\$�L$$�E���C3�;ǉ�$�   �D$ �|$�  �u��d$ �\$�C�<� ���  ���Bx�Ћ؅��  �L$�Q����P|V�҅���   �D$�H�D������\$�L$4� �$�-���ރ��\$�L$D��$�0���L$$Ƅ$�   �0�������Dz�L$$�1��������D{63���|,������L$<�$�������L$,�$�������;�~Ջ|$�L$4�4�Ƅ$�    �j  ��;|$ �|$������L$$Ǆ$�   ������i  �   �L$xd�    Y_^[��]� �L$$Ǆ$�   �����i  3��L$xd�    Y_^[��]� ���SUVW���_3�3���~)�G�<� ��t$�����   �Ѕ�~;�~���;�|�_^��][�_^]3�[���������SW���_3���u�G�D$�����   ���$��_[� ~WV�   3�;�}5�O�<� ��u3��� �D$������$���   �Ѓ���u�^_[� ��t�D$�����$����^_[� ������U����j�h,�d�    P��h  SVW�  3�P��$x  d�    �ً�P4�҃�u,�E�E���$P���\�����$x  d�    Y_^[��]� 3���$�   �|$�����s;���$�  �t$ ~�K�	�3Ƀ�u(;��a  ��E�E���   ���$P�҉D$�A  �;  ��E���   �����$�҅���   �u;�tn�D$TP���4���P�L$@Q��觯��P��$�   �Jg  �E���$V��$�   Ƅ$�  �<� ��u����$��$�   V�#� �L$|Ƅ$�   �bg  ��$�   Ǆ$�  �����Kg  �   ��$x  d�    Y_^[��]� ��$�   R����������#  �L$T�m���L$<�d���L$$�[���C� j j �L$,Q�T$`R�����$�;�����u1��$�   Ǆ$�  ������f  3���$x  d�    Y_^[��]� �L$$�]&������   ��Ph�L$lQ������$�L$TQ��$0  R�����$Ƅ$�  �������$�   �$P��躭����� ����L$$�P�T$(�H�L$,�P�T$0�H�L$4�P�L$l�T$8Ƅ$�   �	f  �L$$��%�����!����   ;�L$������$    �C�<�    ǃ8 ��   ���Rh�D$lP����$�s�����$Ƅ$�  ����������$�   �$P�������L$<�P�T$@�H�L$D�P�T$H�H�L$L�P�L$l�T$PƄ$�   �Ne  �D$TP��$�   Q�L$D���P�T$(R�D$\P��$�   �q�����u�t$ �L$��;ΉL$�&����*����L$ 9L$������E���   ����$�   �$P���҅��D$t�}��t�    ��$�   󥍌$�   Ǆ$�  �����d  �D$��$x  d�    Y_^[��]� ������SVW���_3�3���~:�G�<� ��t,��D$��D$���   ���$P�҅�t��;�|�_^[� 3�_^[� V��N3���u��~7�N�	��t.����   ^��~!��������tj ����������   ^�3�^�������3��yu�I�	��t
����   �������U����j�h|�d�    P��(  SVW�  3�P��$8  d�    ���|$��$�  ������$l  ������$�   ������$�   �����$,  �����$D  �����$�   �����$  �����$�   �|����$�   �p���L$\3��D$ � ���L$4��$@  ����E$;ƋOƄ$@  �L$(�t$$t�0;��  �E�]����D��  �EP��$�   �[����E�E ����t� %�?  �D$��D$    �E�E��������Au�����   �  ~�G�3��T$�t$(RQ���$P��Vj�%d ���}  �؉\$ t9\$u�E ����L$$��D$$    �W�D������ �����@� ��������4� ���@��������A��   �E�E������zt���T��L�������   ���������   �!����������Az~�S;T$(}u�  ����U~�G�3��L$Qj���$PVj�Ic �E�؃��\$ �=�ڍ�����Au,�������Au!�!����������Az��~��]����E������E������Au���D$�����T$|���T$T��T$|�D$   ���T$T�Ʌ���	  ��;\$(��	  �G�D����\$|����A��	  �D$T�����A��	  �O�4�����$�   ��	  ��؋Rh��$�  P���ҋ�L$4�P�T$8�H�L$<�P��$�  �T$@�[`  �G�D��؃��\$�L$l� �$�L#���L$4Q�L$`��'���E��t	�\$L�E�C���L$d�$������L$<�$�P���\$L�E���L$d�$�z�����L$<�$�+���E$�T$D�E0����   ���\$�L$4�E(�$PQ�M��$�   P���\$�D$x�$Q���҄��D$��  �D$4P�L$`�>'���D$t���4  ���L$<�$�������L$d�$���ݔ$$  �E�����E����������������;ݔ$  �D$|���T$l������t�l$T������A��  ����ٍL$\�������L$4�\$,�����|$,����������Au�������'������z������D$D�����D$L������������������;���D$l݄$$  ��������Az��������Au����������D$Tܤ$  ������A��   ������Au����������E0�E$����   ���\$�L$4�E(�$PQ�M��$�   P���\$�$Q���҄��D$tG�D$t���L$<�$�z�����L$d�$�+���D$|������t�D$T������A�  ���D$ �D$ÉD$L��  ;D$(��  �O�����v  �E�L$\�]����z j ����E������Q  �"������j���� �E��������A�-  �]�L$4����zPj �]��� ��\$,�Rh��$�  P����j��Ƅ$D  �5��� ��$�  �\$DƄ$@  ��\  �   �Lj���� ��\$,�Ph��$\  Q����j ��Ƅ$D  ����� ��$\  �\$DƄ$@  �\  ����E�����
�|$l��  ��Ȱ�$����D$,j W��$�   Q��$�  R�����$賗���D$Dj ��W��$�   P��$x  Q�����$荗���}uM��$�   �����4����$�   �$R��$�  P��$�   �S������������   �D$��   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$�   ��$   ��$�   ��$  ��$�   ��$  ��$�   ��$  ��$�   ��$  ��$�   ��$  ��$  ������$  ������$  Q��$�   ����](����z�D$��|$ �  �}$ �  �U$�   ��  �D$,j W��$4  P��$�   Q��$�  R�����$�֖���D$Dj ����P��$L  Q��$�   R��$|  P�����$視���}��   ��$�   ������4����$�   �$Q��$�  R��$�   ������!�����w  ��$,  �����4����$L  �$P��$�  Q��$<  �U�����������  �}$ �D$t	�E$�    �E�L$ �U����{���E��t�T$�R����E ���|$��  ��  ��$�   R��$�   P��$4  Q��$�   R�0& ��$�   P��$  Q��$\  R��$�   P�& �� ��$  Q��$�   �����E(��������A��  �E0��$�   ��$�   ��(�\$ �ă��}�\$0���$�   �H��$   �P��$  �H��$  �P��$�   �H��$�   �ĉ��$�   �H��$�   �P��$�   �H��$�   �P�Hu�\^����E]����@���  �}��   V誜 �����D$,tBS虜 ����t5�E0�t$,���\$�x�E(���$�#���������   ��$�   �|$l��}�΋������&���T$�$������&���T$���$�������:���   �|$ ������D$L�E���|$�D$ ��   ��������}$ �D$������U$�   ������}$ ���D$������M$�   �����}$ �D$������U$�   �����E$���D$�w����    �l����E�E��t����E ��t�L$$��ˉ�����E�|$ uE�E��$�   ;Et4�E0�M$�U���\$�E(�$Qj ��R���\$���$P�����D$����؍L$4Ƅ$@   �V  �L$\Ǆ$@  �����V  �D$��$8  d�    Y_^[��]�0 ��ɪn�e�  �������������U����j�h��d�    P��   SVW�  3�P��$�   d�    ���_3�;��D$F�\$P��  �O��E��������A�  �������  �E��P薔���E�E��;Ɖt$H�t$Lt� %�?  �D$H9w ~�G�3��L$H�EQj���$P��Sj�~W �W���D������� �����@� ��������4� ���@��������Aus�E�������!��������Az��~������U�R���a����������Az@�V;T$P}7�  ���A�U~�G�3��L$HQj���$PSj��V ��������E�U��t9t$Hu����D$L��2�O������A�I  �T������:  V�؋�������؅��<  �L$d����L$TǄ$�       �����Rh�D$tP��Ƅ$�   �ҋ�L$T�P�T$X�H�L$\�P�L$t�T$`�DT  �G�D������\$�L$t� �$�5���L$TQ�L$h�w���E��t���L$l�$������L$\�$�B���E8�M����   ��(�\$ �D$t�E0�\$�E(�\$�E �\$�E�$P���$Q���҈D$F�E��t�L$L��Ή�L$TƄ$�    �S  �L$dǄ$�   �����wS  ���u.�������Dz#�D$F�؊D$F��$�   d�    Y_^[��]�8 �D$P�X�;�u��������D{��E8�]��(�\$ ���E0�\$�E(�\$�E �\$�E�$R���$S�������D$Ft���u���|�;t$P�{����O���E��������u������Z����D�������D�K���V���������V�ϋ������ۋ��,������$�����&���T$���$������&���T$���$�D$W�Q����L$G:�uO�������S�{� V���s� �����������������E8���\$�x�E0�s�$���������������D$F �����E8�U�E��(�\$ ���E0�\$�E(�\$�E �\$�E�$R���$P�Ʋ����$�   d�    Y_^[��]�8 ��������������SUW���_3��������tMV�O�����O�J���3���~(�d$ �O������   �ЋO������;��|܋W�ڍ���^�������_��][��U����j�h�d�    P��   SVW�  3�P��$�   d�    ����P4�w3���3�;�D$X��  ;���  ;E��  �E ;�t����?  �T$D��L$D��9O ~�O�ER�F�uV���$QPj�D$h�`R ������؉\$@t��ua�G�E�\$\�L$\�D���Q���\$� �$V��������t2�  �D$\�U~�G�3��T$LSV���$PRj��Q ���D$@�؋G������  ��Rh�D$tP���ҍL$tǄ$�       ����\$L�L$t�o���\$\�L$tǄ$�   �����O  �D$\���D$L��������D�D  �G�L$@�ȍ��T$l�@�T$d��������Dz��������Dz���������E�   ��������������4��;������Au$���E��������������������Au���V���R�E��������������������������Dz�������$������������Dz�������������Dz�������������u��������������Dz����߃�u�   �E ��t9L$Du����L$H��D$H    �M�}����   �D$HPV�uVQW�����$�ҋЅ҉T$D��   ����   �D$\�d$L�D$d���D$l����������D��   ��������D��   �E���������D$L��|l�\$X3Ƀ�|C�S������F��    �@��� �����X��@����X��@����X��@����X�u؋D$L�T$D;�}����;��L���\��|���Ƀ�u����؋E ��t�L$H��L$@���$�   d�    Y_^[��]� ������������3���$�   d�    Y_^[��]� �Ë�$�   d�    Y_^[��]� ��U�l$��V��~Q�|$ tJ�FS�^W�<(;�~�y���;�}��;�}P����x���T$�F��    Q�NR��R�;� ��n_[^]� ��������������VW�|$����|F�F;�?S�^;�u����;�}P���x���F�F+ǃ�PW�GP����x���T$�N���[_^� ���������VW�|$����|F�F;�?S�^;�u�`?��;�}P���4����F�F+ǃ�PW�GP�������T$�N���[_^� ���������j�h�d�    PQ�  3�P�D$d�    j(�������D$���D$    t���~����L$d�    Y���3��L$d�    Y���������������j�hK�d�    PQVW�  3�P�D$d�    ��j(�t������D$���D$    t���
������3����D$����tW���P����ƋL$d�    Y_^���������������V���(����D$t	V��������^� �̋D$Pj �������� ��������������U��V�u��2Ƀ��  S�\$���  ��5��������D��   �F���W�   |q�{�W�����D��   �G��_�����A��   �����D{k��_�����A{_�W����D{Z�G�����A{N�W����D{I�G�_����A{<���F��� ;�|�;�}.������D{$���\������A{��;�|����������;���u/9u$�}}V�������� |�G    SV������_[^�]� _[^��]� ^��]� ��[^��]� �������U����j�h��d�    P��   SVW�  3�P��$�   d�    �����   ��3�;���  ��P0j���ҋ�Ph�^�L$DQ�Ή|$$�҃���$�   ��   9~�{  �F�;��n  ��Rh�D$TP���ҍD$TP�L$HƄ$�   ����E��u���L$L�$�H������L$\�$�������Bp�����$��;ǉD$ t%�>�L$D��l�����E������ɋ��\$�$�ҍL$TƄ$�    �\H  ��  �EW���T$8�L$P�$�������u=�E���L$L�$�������� ��������Au��$���L$L�$�S����\$,�D$,j���L$P�$�z������1  �F�D$,WW���$P�KQj�I �V���F�����D$H�L$4�э���������z0�L$D��Ǆ$�   �����G  3���$�   d�    Y_^[��]� �Q����t��������D��{�C3�;ÉD$�L$(�L$$��   ���D������\$��$�   � �$�/���D$,���L$|�$Ƅ$�   �����\$4�L$��Rh�D$dP���D$4���L$l�$Ƅ$�   �%����L$����   �T$$R�T$,R���$�Ѕ��D$ u1��$�\$4����z��;�}�N���T$��D$    �l$�L$dƄ$�   �mF  �L$tƄ$�    �\F  �D$3�;�u�T$�T$$�L$�D$    �
9L$ ��  ;���  �V��P�L$X�z����D$��P�L$8Ƅ$�   葛���L$$Q�L$XƄ$�   �+����T$,R�L$8��A���F�D�+�P���S�L$\�����F��    �L$�LQS�L$<�����F�\$<PW�L$\�w����FPW�L$<�y����|$( t�T$(R�L$X贓���FD$�L$4P�A���L$,Q�L$8�uA���L$D�L���;\$<}�D$8�؃����\��;\$<|�F�؋N��    Rj Q�x� �N���y |�A    �D$X�T$\PR������F�@�N�T$4R�ЋL$��t	��Bj�ЍL$4Ƅ$�   �����L$TƄ$�    �C�����D$    �>�L$D��l�����E������ɋ��\$�$�ҍL$DǄ$�   �����pD  �D$ ��$�   d�    Y_^[��]� ����U����j�h�d�    P��   SVW�  3�P��$�   d�    �ى\$$�L$d�/���3��L$T��$�   �����u;�Ƅ$�   �|$ t9~|�~�}3�;�t9O|�O�C���D$0��   �C9t�����   WV�҉D$ 3�;��m  9L$ �c  �C�@���\$�L$t� �$����C���Rh�D$DP�ҋ�L$T�P�T$X�H�L$\�P�L$D�T$`�DC  �D$TP�L$h�
������  3�9w��  �����O��<���L$\�$�������L$l�$�G�����U��;r|��  ��  �D$D�$�L$H�L$L�L$P�D$4%�L$8�L$<�L$@3�;�Ƅ$�   ��  ������D$4#��E����L$D#��t$(�D$,����D$,3�9L$P|�L$L9L$@|�L$<�T$$�J���VP���   �Ѓ��(  D$ ��t�l$ ����   �L$$�Q�D��ڃ��\$�L$t� �$����D$$�H����Rh�D$tP�ҋ�L$T�P�T$X�H�L$\�P�L$t�T$`��A  �D$TP�L$h�'	����tB3�9t$<~6�L$8��<���L$\�$�2������L$l�$��������;t$<|͋}�t$(�G��~����P�B���ЋL$8�T$<QR���L����M��t$�A��~����P�B�ЋM�T$H�D$LRP�����;\$0������u�#�E3�;�t9H|�H;�t9O|�O�L$ ���L$$����   ��3���tK;�tG�F��~?;�~�N�3�;�~�@�F�D���3����Q�P�Q�P�Q�P�Q�P�I�H9|$@Ƅ$�   �D$4%t �D$8;�tWP�L$<�%�|$8�|$@�|$<9|$PƄ$�   �D$D�$t �D$H;�tWP�L$L��$�|$H�|$P�|$L�L$TƄ$�    � @  �L$dǄ$�   �����@  �D$ ��$�   d�    Y_^[��]� U������$SVW�}����^�D$    ��  ;���  �M����  ;���  �D$P�T$R��s������  �EPW�N�D$   �����;���   ��u(�L$��Q���;���T$R���~;���D$_^[��]� �F�����D$��������Dz&�ٍL$ ��Q�D$�N�\$$�A;���D$_^[��]� �l$�L$ Q�N���\$$�;���D$_^[��]� ��uF�V����D$��������Dz
�����D$��l$���D$ �\$ Pj �N�c����D$_^[��]� �N�����D$��������Dz���D$��l$���T$ �T$ ��R�GP�N�\$0�����D$(�v�O�{��+у���|<��+у������D����@��� �����X����@��X��@����X��@����X�u�;��΃�;����\��~��؋D$_^[��]� ��������������U����j�hz�d�    P���   SVW�  3�P��$�   d�    ��F ���^�\$(�'  �K;��  �}����������
  ��Rh��$�   P���ҍ�$�   Ǆ$       ��������  ��O�W�D$<�G�L$@�T$D�D$H��$�   Q�L$@Ƅ$  �8�����L$<�v  �W������L$<�e  ��$�   R������N  �D$<�L$@�T$D�D$l�D$H�L$p�T$t�D$xj �L$@Ƅ$  �D$$�����D$���������� j�L$$Q�����$�m�����t!�D$ ��|;��Vj �L$p�<�������j�L$@����� j�L$Q�����$�'�����t&�D$��|;��Vj�L$p�<��V������l$�L$l�d������a  �L$ ���U  �D$;��I  ;��A  ����p����$�   P�L$p�����t}�~j �L$@������ ��N�4�j�L$@������ ��L$lƄ$   �;  �L$<Ƅ$    �;  ��$�   Ǆ$   �����p;  �   ��$�   d�    Y_^[��]� 3�9|$ ~&�V����t	��Pj�ҋF��    ��;|$ |ڋ|$�_;\$(}*�N����t	��Bj�ЋN��    ��;\$(|ڋ|$�W�^R���p-���G�NP�d-���|$  ��   +|$ ��$�   ��W�����L$+L$ Ƅ$   ��Q��$�   �%����L$ �F���D$+�R��P��$�   Ƅ$  �L����L$ �F�ȋD$+�R��P��$�   �;������{���{ |�C    ��$�   ��$�   QR��� ����F�@�N��$�   R�ЋD$+D$ ��$�   �D$�D$     Ƅ$   �%�����$�   Ƅ$   �a����~j �L$p������ �����At*�|$ u�~j�L$p�������������At�D$' ��D$'�D$;D$ ~"�N�|�j�L$p�������D$����At�D$ �L$,�o����L$|Ƅ$   �^����L$\Ƅ$   �M����L$LƄ$   �<����|$' Ƅ$   �S  �~ ~�V�:����$�   ��   �L$LƄ$   ��8  �L$\Ƅ$   ��8  �L$|Ƅ$   �8  �L$,Ƅ$   �8  �L$lƄ$   �8  �L$<Ƅ$    �8  ��$�   Ǆ$   �����r8  3���$�   d�    Y_^[��]� ��Ph��$�   Q���ҋ�L$\�P�T$`�H�L$d�P��$�   �T$h� 8  �L$\�g������ ���j ��$�   P���>�����L$L�P�T$P�H�L$T�P��$�   �T$X��7  �L$L������������L$P�D$L�T$T�L$0�L$l�D$,�D$XQ�L$0�T$8�D$<������������|$ ~-j�L$0����j�L$P�D$,����� �T$(�����D�m����L$,�������\����D$LP�L$`��������   j �L$0�Z���j ��$�   ���J�������L$T�$�D$0�������L$d�$�F����L$(�j�L$0����j��$�   ����������L$T�$�D$0�P������L$d�$�����T$(�L$|��������u<j �L$0������L$L�v�L$,�T$0�D$4�L$|�L$8��$�   ��$�   ��$�   ���$�   �T$\R��$�   ��������   ����   �L$|Q���҅�j ��  ��$�   �K����L$\� ���$�����<�����
����|$ ������F���t	��Bj�ЋN�    �V�B�Nj �Ћ�Bj ���Ѓl$�|$ �7  �L$�F�Q;������Q��豰�����D$(�������Rh��$�   Q���ҋ�L$\�P�T$`�H�L$d�P��$�   �T$h�M5  �L$\�������M����D$P��$�   Q���h�����T$L�H�L$P�P�T$T�@��$�   �D$X�5  �L$L�H����������N�T$�<�j�L$p����� ���\$��$�   ��$�������L$,�P�T$0�H�L$4�P��$�   �T$8�4  �L$,������������j �L$`����j ��$�   ���������D$LP�L$`������j�L$0��   �y���j��$�   ���i�������L$T�$��$�   �������L$d�$�b�����$�   ��L$|�P�������   j�L$0����� ���L$T�$�l�����'����A������D$��������V������   ��Pj����   �~�L$p������ ��L$��������~ �����8L$������~����   ����j��$�   ���������|$ ��   �D$|P�L$`��������   �L$(����   �D$|P�҅���   j��$�   �5���� ���L$d�$������'����A������D$��������N����t��Bj�ЋD$�N��    �F �V�R�N��P�ҋK��P��Q���҃l$��F �N�|��j�L$p����� ��~j �L$@����� ��F �Vj�L$@�|���}���� ����2g���L$LƄ$   �12  �L$\Ƅ$   � 2  �L$|Ƅ$   �2  �L$,Ƅ$   ��1  �P������������U����j�h �d�    P���   SVW�  3�P��$�   d�    ���Ph��$�   Q���ҋE�8��Ǆ$       thPf���G����t�߉�$�   �	3ۉ�$�   �M�9��thPf���nG����u3��ۉ�$�   t;ދ�t�2�����+f����t;���t������f���U�: t���  �E�8 t���  �Ej����$�   �$�~�������  ;�t;��D$\   u�D$\    ��4���$�F�EPj�L$@Q�����$�����؄ۋD$0t����  ;F��  P��$�   R��輫���D$0��Ƅ$   �U  ;F�L  �N�<����>  ��Rh��$�   P���҄�Ƅ$   ��$�   tj �V���� �8��$�   P������E��u$����$�   �$��������$�   �$�:���3��T$4�ۉ�$�   ��$�   �   j����$�   �$�J�������   ��D$4���   ��$�   P��$�   Q�����$�҅���   �D$4����$�   �$�������'��$�   ����Az3�W����� �\$4�   �D$4���$������<��$�   ������   Ƅ$   �/  ��$�   Ƅ$    ��.  ��$�   Ǆ$   ������.  3���$�   d�    Y_^[��]� ����$����$�   �$�����\$4��$�   ����uj �j������ �\$43���D�D$`�|$d�|$h�|$l�D$<�|$@�|$D�|$H�%�D$p�|$t�|$x�|$|�D$L�|$P�|$T�|$X9�$�   Ƅ$   ��  9�$�   ��  �D$0��;�~
P�L$d�Z���F+D$09D$H}
P�L$@�Z���D$h��9D$|}
P�L$t������D$D��9D$X}
P�L$P������\$\;�u!�F�L$0��;�t	��Bj�ЋN�T$0�<��|$0 ~F��t�F���������L$4�D$4Q��V��P�L$d�{���N��R�L$t�|)����;|$0|���$�   P�L$d�{���N�T$0��P�L$t�N)���MQ�L$t�A)����$�   R�L$@�P{���EP�L$P�#)���|$0��;~}K��$    ��t�N����?���T$4�D$4R��F��Q�L$@�{���V��P�L$P��(����;~|��F�N��R��  j��$�   ����� �\$4����Dz�D$0W��$�   ����� �\$4����Dz9|$0t$j��$�   ����� �\$4����D�D$0zU;FuP�L$LƄ$   �h����L$pƄ$   �W����L$<Ƅ$   �|���L$`Ƅ$   �|����$�   �����9D$l}
P�L$d��W���F+D$09D$H}
P�L$@��W���D$h��9D$|}
P�L$t�����D$D��9D$X}
P�L$P�����|$0 �\$\~F��t�F����������L$4�D$4Q��V��P�L$d�y���N��R�L$t�l'����;|$0|��EP�L$t�V'���|$0;~}P��t�N����|����T$4�D$4R��F��Q�L$@�Ay��;|$0u�UR��F��Q�L$P�'����;~|��F�V��P�L$P��&����$�    u4j(��s�����D$4��Ƅ$   t	���o����3�Ƅ$   ��$�   ��$�   ��u/j(�s�����D$4��Ƅ$   t	���0����3�Ƅ$   �؃|$\ u^�N��t�F��~��    Rj Q荳 ���N�ɍ~t�G��~���Pj Q�j� ���~ |�F    � |�G    �L$d�T$h��$�   QR�N�����D$t�L$xPQ�N貮���T$@�D$DRP�K�����L$P�T$TQR�K莮���E�M�03�9t$X�%�Ƅ$   �|$Lt �D$P;�tVP�L$T�%�t$P�t$X�t$T9t$|Ƅ$   �|$pt �D$t;�tVP�L$x�%�t$t�t$|�t$x9t$H��DƄ$   �|$<t �D$@;�tVP�L$D��D�t$@�t$H�t$D9t$lƄ$   �|$`t �D$d;�tVP�L$h��D�t$d�t$l�t$h��$�   Ƅ$   �(  ��$�   Ƅ$    �(  ��$�   Ǆ$   �����(  �   ��$�   d�    Y_^[��]� ����j�hP�d�    P��DSUVW�  3�P�D$Xd�    �|$h�_3�V�L$p�t$d�\$�N���� ��\$ �Ph�L$(Q����;��D$`�Q  ��$�   V�D$<P���)���j���D$d����� �L$8�\$�D$`��'  �D$���L$0�$�D������L$t�$������\$����   ;w��   �O�,���l$h��   hPf���=����t}�D$���\$�L$X�D$0�$�c����T$|SR����̉�P�Q�P�@�QU�D$|�A��������L$H�D$`�'  ;w}
�O��    �U �Bj�����8�D$h    �L$Q��$�   � #���T$hR���u����|;w}
�G��    �D$��;t$�\$ ������L$(�D$` �&  �L$l�D$`�����&  �L$Xd�    Y_^][��P����������U����j�h��d�    P��   SUVW�  3�P��$�   d�    �ًs3��kU�L$h�D$S �t$T�D$h%�|$l�|$p�|$t�%��S�L$X��$�   �D$X�D�|$\�|$`�|$d��D�   9EƄ$�   |�E9{|�{;���   �D$X�4�����   hPf���;����tr�D$h�D����\$��$�   ���D$_�$�����SU���̉�P�Q�P�@�QVƄ$�   �A��������L$tƄ$�   �9%  ��Bj������L$h�T�R���<!���D$X��Q���Ms����;|$P�C���3�9|$`Ƅ$�    �D$T�Dt �D$X;�tWP�L$\��D�|$X�|$`�|$\9|$pǄ$�   �����D$d%t�D$h;�tWP�L$l�%�D$O��$�   d�    Y_^][��]�U����j�hΪd�    P��   SVW�  3�P��$�   d�    �ٍK�u���s3�9~t�F;�t�WP�B���Љ~�~�~�L$XQ�M�T$TR�|$X�|$`��o����;���  �M�D$P�|$�|$X�|$P��X������ty�L$TQ�M��X������te�M�T$LR��X������tQ��$�   �#  �M��$�   PǄ$�       �Y����$�   ��Ǆ$�   �����q#  ��t�MV�`�����D$3�����   ���  �L$0Q�M�D$4    �f:������tS�T$0R��V�������D$$t�D$$P�K�Nq���/h4<h <h�  h�;�����L$@����t	��Bj��3��D$��;��{�������  �K���h  ;��`  �K ��;��R  �L$<�����   �L$��$�   �����{ Ƅ$�   ~�K�	�3ɋ�Rh�D$dP�ҋ�L$�P�T$�H�L$�P�L$d�T$ �@"  �L$�7����D$���?  ���C���L$�T$�\$$�D$�L$<�\$d�L$ �T$@�D$D�L$H|;s}�S���3ɋ�@h�T$tR�Ћ�L$�P�T$�H�L$�P�L$t�T$ �!  �L$�����\$\j�L$@������ �T$4�D$$������D��   j �L$����� �\$4����Dzpj �L$@����� �\$$����zXj�L$����� �D$$��������z:�D$\�D$d������A{�����D$4����������4������u�C�����
���D$\��ًD$��;��������4�Kj�\$h���L$�\$(������ �T$4�D$$������D{Aj �L$������ �D$$��������Au#�D$4���������\$d����Az�S�D$����؍L$Ƅ$�   �g   �L$<Ǆ$�   �����S   �M��  =�e�}��������ǋ�$�   d�    Y_^[��]� ���V���U���L$�FQP������^� ����j�h��d�    P��SUVW�  3�P�D$d�    �ًkj(�l$��h�����D$3�;Ɖt$$tU���������3�S���D$(������;����~:��|/;s}*�C����t ��Bd�Ћϋ��cT���OUQ���w����l$��;�|�;ou�{  ~�[�3�S�������ǋL$d�    Y_^][���������������V�t$��thHg���5����t��^�3�^���������������̸Hg�����������j�h(�d�    PQVW�  3�P�D$d�    ��t$�b2����<�`/�F�d/�N�h/�V�l/�F�`/�N�d/�V�h/�F �l/3��N$j�N0�|$�~(�4_�����   ���   �ƋL$d�    Y_^������́�   VW�y0��$�   W�D$P�3`����    �_�   ^�Ā   � ����������SV�t$��;�t5WV�>���F(��0���{0�    �C(�_t���C(��u^�C(   [� ��^[� ��������V���   ����<tT�F3҅�tK��    ;�t�Ћ��   ��u�^��8����t���   ���   �	���   �Vǀ�       ǀ�       ^�8�������j�hX�d�    PVW�  3�P�D$d�    ���t$hp=V��d�������Cd��V���K4���L$��a����P4�L$Q���D$    �ҍL$�b����thd=�L$ ��i���L$�c��PhH=V�ld��h4=V�ad�����GP���j��h�&V�Hd���O(Qh=V�9d����B8�����Ѕ��=u�=Ph�<V�d��������c���L$�D$�����H`���L$d�    Y_^��� �����+3���   �����̃� VW��~h`/W��{������u �D$,��tht>P�c����_3�^�� � �D$P�Hg�%/��PW�n|������u �D$,��t�h(>P�dc����_3�^�� � ��B8���Ѕ�tU�L$Q�Hg��.��P��T$R����ҋ���.��P�|������u$�D$,���o���h�=P�c����_3�^�� � _�   ^�� � �������̋��   ���������̋��   ���������̃�V�����=0hu���   ��L$Q���9.���L$���P�Q�P�@�Q�A��^��� �����̋���3�=0h�����������������̸0h�����������V��������>�`/���   �d/���   �h/���   �l/���   3����   ���   ���   ���   ��^�������VW�|$��;��Y  ���   S3�;É��   tP�g}�������   W�������9^(�G�F�O�N�W�V�G�F�O�N�W�V�G �F �O$�N$��   9��   ��   9��   tx���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   QR�� ���   ���   �����   ���   [_���   ��^� �`/�V�d/�F�h/�N�l/�V�`/���   �d/���   �h/���   �l/���   ���   ���   ���   ���   [_��^� V���/�����   �   �D ^�������̋L$h�>�be���   � ���������̃��  3ĉD$�D$VP���E�����tS3�9��   ����tD3�9��   ����t5�Ƹ   h`/V��w������t�D$P�0h�l+���L$QV��w�����L$3҅���^3̋�蓜 ��� ���V�t$WV���������_��h`?V�_�������   P����e��h�&V�d_�����   Qh<?V�R_�������_��_^� ��̸   ����������̋��   ���   PQ�L$�C����� ���V���   ���   WPQ��z���|$���ω��   �e&�����   ���   ���   RP���jB��_��^� ��j�h��d�    PQVW�  3�P�D$d�    ��t$j�0H���|$ �|?���   P���D$    �P+�����   ���@  ���   ���@  ǆ�@      �ƋL$d�    Y_^��� ���������|?�H������̋��@  ����������V�t$2���}����9��@  r���@  �;��@  s���@  �^� ������������̋T$2�;��@  s3�;��#��@  �� ��������������̋��@  ;��@  ���V�񋆘@  ���@  3�;�Wv+��Ћ|$;�v����v���@  ��L$WPQ��� ����@  ��_^� ����V���()���D$P���\*�����$�������^� ����������̀|$ VW�|$��u����(��V���"*������(�����d$�����_��^� ���������j�h��d�    PQV�  3�P�D$d�    ��t$��Y���N�D$    ��Y���ƋL$d�    Y^���j�h�d�    PQV�  3�P�D$d�    ��t$�N�D$    �X�����D$�����X���L$d�    Y^�����������V�t$Wj j��h � @���������u_^� SW����]���؄�t��W����]���؋�������u2ۊ�[_^� �������������̃�UVW���SX���n���IX���|$3��D$�D$�D$P�L$Qh � @���5�����u	_^]��� �|$S�Ä�tV���M���؄�t
U���M���؋�������u2ۊ�[_^]��� ����������V�t$��thi���[)����t��^�3�^���������������̸i�����������V�t$��th j���)����t��^�3�^���������������̸ j����������̋L$j�V����� ��������������̃�SV�t$�D$P���D$ ��E���؄�tV�D$�Ȁ���wH<u93��T$�D$�D$R�D$Ph � @��������t �|$����������u2�^��[��� ^3�[��� V�������D$t	V�K]������^� ��j�h�d�    PQ�  3�P�D$d�    h�   �[�����D$���D$    t���k����L$d�    Y���3��L$d�    Y������������V�t$��th0h���'����t��^�3�^����������������j�hK�d�    PQVW�  3�P�D$d�    ��h�   �qZ�����D$���D$    t����������3����D$����tW�������ƋL$d�    Y_^������������VW�|$��t5h0h����&����t%�t$��th0h����&����tW������_�^�_2�^�������������V���   ����>t	P�t������������D$t	V�[������^� �������V���|?��B���D$t	V�u[������^� ������������j�h{�d�    P��@  ��� �  3ĉ�$�@  SVW�  3�P��$�@  d�    ���P3�W�҅���   ���   ���   ���ĉ���   �P���   �H�P�����;���   ���_����;�tshHg���%����u��Pj��3��ҋ��TV�L$�����F(��R$��$�@  �C(��0�{0�    �D$�P���ҍL$Ǆ$�@  �����D$|?�A������ǋ�$�@  d�    Y_^[��$�@  3��Γ �Ĵ@  �������������̋��   �L$Ph�?Q�
]�����   � ���������������SVW����%�����   �����   ����   t���   ����H�S�����Cu�_^��[��������������̋D$SU�ً��   V3���~9W���$    ����   �<�    �P�T�����   �P����S����;�|�_^][� ������������QS�\$UV���   WUh@S�t$��U�������EU��3���~U��t$���   �4����IT����u��7Ph�?S�U�����N�)T����u��7Ph�?S�tU������;�|����#U��_^][Y� �����������QU�l$Vj ��jh � @�͉t$�������u^3�]Y� SW���   W���WS���؄�t&3���~ ��t�D$���   ��U�������;���|����~����u2�_��[^]Y� ���j�h��d�    PQV�  3�P�D$d�    j��U�������t$3�;��D$t���m ����?�ƋL$d�    Y^�������j�h�d�    PQVW�  3�P�D$d�    ��j�U�������t$���D$    t��� ����?�3����D$����tW���-���ƋL$d�    Y_^���������VW�|$��t5h j���"����t%�t$��th j���"����tW����,��_�^�_2�^�������������V����?�B'���D$t	V��V������^� �����������̃�V�D$��P�i����P���������t%hi���!�����D$t��RP����^��� �D$^��� �������������S�\$��V��~[U�l$��|QW�|$��|G;�tC�F�+;�9;�5�N�;�~�;�}��P���6����F��    R��Q��R辔 ��_]^[� ����SV�t$��;�tn�FU3�;��k]^��[� 9C}P����9kt�F;ŉC~�W����t$�v�{��    ��V���3V����V�O�'V����;k|�_]^��[� ^��[� ���������������VW�|$����|`;~}[�NS��    ��m����F�3ɉ�H�F+ǃ�P�OQW�������V�N�L��3���A�V�F�L��Q���y/���F�[_^� ���������������SU�l$��;�t0VWU�*���E(���u0�{0�    �C(�_^t���C(u�C(   �Ÿ   U���   ����]��[� �����������VW�|$��t5hi���Z����t%�t$��thi���B����tW���f���_�^�_2�^�������������j�h&�d�    P��V�  3�P�D$d�    ��t$����3��@�D$$ǆ�   h����   ���   ���   �D$P�i�D$(�����N�P�V�H�N�P�V��/�F��/�N��/�V ��/�F$�F(   �ƋL$d�    Y^�� ���j�hX�d�    PQV�  3�P�D$d�    ��t$�@���   �D$    �������D$�����`����L$d�    Y^������������������V��F�V;�uN��    ��   v��|�  ;�}�������   ��;�}5P���օ���N�F�ȃ��N^ËV��������N�F��R���	-���N�F�ȃ��N^���������j�h��d�    PQ�  3�P�D$d�    h�   �EP�����D$���D$    t��������L$d�    Y���3��L$d�    Y������������j�h��d�    PQVW�  3�P�D$d�    ��h�   ��O�����D$���D$    t���������3����D$����tW�������ƋL$d�    Y_^������������V�������D$t	V�kQ������^� �̃�UVW�|$��D$P�L$Q3�h � @�ωl$�l$蔅����u_^3�]��� �|$S�Ä�tV�T$R�ωl$ ��:���؄�t@9l$~:�Ƹ   ��    W���������������؄�t��;l$|���F��P���b������+y����u2���[_^]��� ���������K� ������������K� ����������̃�`�  3ĉD$\�D$pU�l$h�D$�D$l��W�|$t�l$�2  SV�����������݃�@�t$$�D$�\$ vW�Hh�����D$��L$,�L$����I ��Wt�������RP�t$0�F� ���#SP�:� WUS�2� ���l$��   +߉\$ ����l$�\6;\$w_����t$;\$s�7PV�D$0�T$$����}�t$(���D$VP�T$$����}WVU�ȑ ����\��\$��;\$v��t$$�L$WQU蠑 �l$$�\$,�D$���,����t$WVU耑 ����@v	V�g����^[�L$d_]3�誈 ��`�������������U�l$W��;���   �M�    S+�V�_�D$��D$Ù����������M|F��������z����Q�����z����Q�����z����Q�����z��� ;�~�;�w������z���;�v�����G��;���_�q���^[_]��������U�������   ��SVW��  ���  �D$    �؍|���\$��+�������w)S����������D$���D$�B  �\�����   �����Í������z����������z����������z�����Ӌ��I ;�v��;�s������t�;�w��;�w������t��;�v������{�;�r;�����u���뮃�;�s��;�v������D{�;�r��;�v������D{��+L$��+�����;�|-�D$;�s�L$�D�����   ���L$;������������;�s�D$�T�����   ���D$�\$;������������_^[��]�����������Q����   ���   SUV�؍p�����D$��t	�D�������� ��tQ���D$�L;΍,�w:;΍�s��Z����z���������z��L	�] ����N;�vʋD$�] �^�][Y�������������̃|$ u�D$W�|$�K���_ËL$�D$������������������V���T$�\$�����$覹������T$�\$�N�0'�$船����^����̋��L$���Q�P�Q�P�Q�P�Q�P�I�H�L$��P�Q�P�Q�P �Q�P$�Q�P(�I�H,� ������������������������������VW���׺���~���ͺ������0'�_^��������������̋D$���Q�P�Q�P�Q�P�Q�I�P�H� �������U������SVW��3��;�����tf�L$�η���]3҅�t�F���3ɍÅ�t�F ��F�F���ʃ����0�����P����X��F(���P����X��X�|Ń��؃�|�3���_^��[��]� �|$ �T$����tI��A��   �A�����Au~�B�Y����Auq�A �Z����Aud�B�Y����AuW�A(�Z����A�C��uE�A�����u9�B�Y����u,�A �Z����u�B�Y����u�A(�Z����u�� 2�� ������̃�SV��2���������   U�l$����   W�|$ ����   ;���   U������� W�\$������U�΋������W���������D$���U������� W�\$���ٻ��U�΋��ϻ���W����û���D$_�]^�[��� ^��[��� ]^��[��� ��_]^[��� VW���7�������   �|$���$�����tz������z���F�_����z�G�^�F�_����z�G�^�F�_����Au�G�^�F �_ ����Au�G �^ �F(�_(����Au/�G(���^(����_^� ���Ϸ���~���ŷ������0'�������_^� �������������SV���g������t$����   �T�������   ������Au���C�^����Au�F�[�C�^����Au�F�[�C�^����z�F�[�C �^ ����z�F �[ �C(�^(����zO�F(���[(�����^[� �������tW�   ���_������^[� ���۶���s���Ѷ������0'�������^[� ���������SV�t$��W���p�������   �|$���]�������   ������Az�����G�^����Az�F��G�[�G�^����Az�F��G�[�G�^����u�F��G�[�G �^ ����u�F ��G �[ �G(�^(����u�F(���[(�ȿ��_^[� �G(���[(赿��_^[� ���ص���s���ε��������0'�苿��_^[� �����U����j�h�d�    P��hSVW�  3�P�D$xd�    �ى\$��D$ 3���I �\$���  �{V���Y������$V���K������L$D�$�\����]��V��Ǆ$�       �#����M���$V�������L$4�$�%���j �D$(P�L$<Ƅ$�   �m����} �D$tR�|$ uK�MV�ӷ���\$�L$V�ŷ���\$����{$V��買���\$V��覷���\$�D$ ����Au�D$�L$$Ƅ$�    �����L$4Ǆ$�   �����|����D$����������} t$��t�|$ t��L$xd�    Y_^[��]� 2��L$xd�    Y_^[��]� ������������̃|$ V����   �ͽ����tx�L$�������Au���^����Au��^�F�Y���A��Au�^��^ ����Au�A�^ �F�Y���A��Au	�^�^� �^(����AuU�A��^(^� �D$���P�V�H�N�P�V�H�N�P�V��N�P�V�H�N �P�V$�H�N(�P�V,�^� ��U������tS�] ��VW�}�D$' t���޼����u3ۋ������w�����������0'��E��t�   �E�}����  �M����  �u����  ��t�9M�{  �L$P��������T$�T$�L$P�$蹰���M$��t����$�>����t�E$    �]���\$,~�E   �} �D$'��   ����U|S������Dz~��    ����D$' ����DzY����D$' ����DzM����D$' ����DzA�����D$' ���~������Dz'�����4��D$' ���2�_^[��]Ã�����������~�E���P�D$,�D$TVP�� ���} t!���4��D$P���\$P�D$X���\$X�L$`�\$`�E$��t
P�L$T�ܬ���]�L$P�T$T�D$X��ۉL$h�L$\�T$l�T$`�D$p�D$d�����L$t�T$x�D$|��  �} �.  �}$ �4  ���L$,�΃��T$0��$����Dz
�D$' �   �T$(R�D$<VP�K� ���t$<�M$��Q�L$<�D$<���\$<�D$D���\$D�L$L�\$L�����D$8�T$P����z�\$P��T$h����Au�\$h����D$@�T$X����z�\$X��T$p����Au�\$p����D$H�T$`����z�\$`��T$x����Au�\$x����������}��  �uV�L$T� �����V��L$l����������|܍L$PQ�M�9����D$'_^[��]ËT$,�փ��T$0��$����Dz
�D$' �   �D$(P�L$<VQ�� ���t$<���D$8���T$8�D$@���T$@�D$H�����T$H���T$P����z�\$P��T$h����Au�\$h������T$X����z�\$X��T$p����Au�\$p����T$`����z�\$`��T$x����Au�\$x������(����L$PQ�M�I����D$'_^[��]Ã}$ ��   �d$ �T$(R�D$<VP���=� �M$��Q�L$<�-����D$8�T$P����z�\$P��T$h����Au�\$h����D$@�T$X����z�\$X��T$p����Au�\$p����D$H�T$`����z�\$`��T$x����Au�\$x������[����}��   �uV�L$T�4�����V��L$l�&���������|܍L$PQ�M�M����D$'_^[��]Ë��T$(R�D$<VP���M� �D$D�T$\������z�\$P��T$h����Au�\$h����D$@�T$X����z�\$X��T$p����Au�\$p����D$H�T$`����z�\$`��T$x����Au�\$x������h����L$PQ�M�����D$'_^[��]Å�t���D$'�D$'_^[��]����������̃��D$S�\$,UV3Ƀ�W�|$<�D$ |v��s�W+$    �|$@ ��   �B��^������u  ��*�����e  �B�^������T  �B�����z�D$@    �D$$���x��� �� ;�|�;�}7�D$<�l$$�|$@���+��d$ ��t��2����z3�����;�|�|$@�|$,���J  �D$(��t�   �t$4����  �L$$����  ���T$0t�,;���  ���D$��  ����|b�,�    �.����D��   ��    ��.�D$ ����Dzx��.�D$ ����Dzl��.�D$ ����Dz`�����D$ ��L$$���  �,�    �.����Dz7�����4��D$ �D$��_^][����D$@    ����������������  �|$@ ��u6�ًD$$�4.SV���$P�m� �L$PUSQ�} ��T$P��� �ɍ4փ����l  ��    �D$��|$,�L$$���΋l$<���|$,����Dz
�D$ �'  ��3҃��4���   ��+ÉD$�}��+�+D$<�K�D$�����Q�����z�Y���W�����Au�_���؋D$��������z���)����Au�)��؋D$�8���Q����z�Y������Au�����D����Q����z�Y��W����Au�_��؋D$$������� �� ;��O���;T$$}D�l$<�|$$��+�+��+��D$����������z���)����Au�)��؃���u���t$�|$, ��������؊D$_^][��Ã|$@ u-�����UVS��{ �L$HUSQ��{ �T$H�����4։|$,��t���    �D$�	��I �\$8�l$,�D$<3҃|$$��   ��+�l$��K+�ލx+����Q�����z�Y���W�����Au�_���؋D$������z���)����Au�)����;�Q����z�Y������Au�����D��Q����z�Y��W����Au�_��؋D$$������� �� ;��[���;T$$}@�D$8�l$<�|$$��+�+��+�������z���)����Au�)��؃���u�t$�|$, ������D$_^][��Ã|$@ �i���_^�D$�D$][����������������̃��D$S�\$0UV3Ƀ�W�|$@�D$ |~��s�W+$    �|$D ��   �F��B��������y  �*��������g  �F��B�������T  ��B������z�D$D    �D$(���x�����;�|�;�}5�D$@�l$D�|$(���+���t�2�������z3����;�|�l$D�|$0����  �D$,��t�   �t$8����  �L$(����  ���T$4t�,;���  ���D$��  ����|b�,�    �.����D��   ��    ��.�D$ ����Dzx��.�D$ ����Dzl��.�D$ ����Dz`�����D$ ��L$(���U  �,�    �.����Dz7�����4��D$ �D$��_^][����D$D    ���������������  �|$D ��u<�ًD$(�4.SVQ�\$<�D$<�$P聱 �L$PUSQ�%x ��T$P����ɍ4�������  ��    �D$��|$0�D$(�����0���|$0����D�w  �D$(��3҃����	  �D$@��+�l$��x��+�+D$@�K�D$ �����\$�A��D$��������z�Y���G�������z�_���؋D$����\$��D$��������z���)������z�)��؋D$ �8���\$�A�D$��������z�Y��������z�����D����\$�A�D$��������z�Y��G������z�_��؋D$(���������;�����;T$(}R�l$@�|$(��+�+��+��D$���
���\$��D$��������z���)������z�)��؃���u���t$�|$0 �W������؊D$_^][��Ã|$D u+����UVS�/v �L$LUSQ�#v �T$L�����4��|$0��t���    �D$���\$<�l$0�D$@3҃|$(��   ��+�l$��K+�ލx+����\$�A��D$��������z�Y���G�������z�_���؋D$��\$��D$��������z���)������z�)����;�\$�A�D$��������z�Y��������z�����D��\$�A�D$��������z�Y��G������z�_��؋D$(���������;��#���;T$(}T�D$<�l$@�|$(��+�+��+���    ��\$��D$��������z���)������z�)��؃���u�t$�|$0 ������D$_^][��Ã|$D �#���_^�D$�D$][�����S�\$(UV3Ƀ|$W�|$8|h�l$0�u�S+����   �B��^�������   ��*������   �B�^�������   �B�����z3��D$������� �� ;�|�;L$}+�t$0��+�d$ ��t��2����z3�����;L$|����3�9t$�D$8~i�l$,�\$(���$    �L$4�T$0���D$$WQR�T$,�L� �D$$Q�L$$SRPQ������� ��t#���   u�D$8�;t$|��D$8_^][�3��2�_^][���̋T$3�9D$j ��P�D$Q�L$ Q�L$R�T$PQR�U����� � ��������������́��   SVW�ٍt$�   ���ŝ������y�$�   �N��t�F�@���Pj Q�n ���L$Q���F    �����؄�tK�FU�n�x;�~���Y}��;�}��;�}P���|���F�Nh�   �T$R�@��R�Kr ���F]_^��[���   � �����j�h�d�    P��SV�  3�P�D$d�    ��L$������D$P���D$(    ������؄�t=�L$,Q�L$�8����؄�t)�D$3Ʌ���j j V��#L$QjPj j������� �؃|$ �D$$�����D$�$t�D$��tj P�L$��$�ËL$d�    Y^[��� �������V�t$��thHk���������t��^�3�^���������������̸Hk�����������VW�|$W���������   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ݇�   _ݞ�   ��^� �����������Q�`/V�񉆸   �d/���   �h/���   �l/j �L$���   ǆ�       ������'�L$ݞ�   ���   ^Y�������(��������SV�t$Wj j��h � @���7����؄�tf���   P���*���؄�tR���   Q����R���؄�t=���   R���z(���؄�t)���   P���*���؄�t݇�   �����$��)���؋��4S����u	_^��[� _^��[� �������������̃�SV�t$W���D$P�L$Q�   h � @�Ή\$�D$    �]a����u_^3�[��� 9\$u�   R�������؄�tL���   P���%���؄�t8���   Q������؄�t$���   R���.���؄�t���   W���
���؋���T����u2�_^��[��� ��������������̋D$h�AP�Q/�����   � �����̸0l�����������VW�|$W���������   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ݇�   ���   ݞ�   ����   �P���   �H���   �P���   �H���   �P_���   ��^� �����������̡`/�艁�   �d/���   �h/���   �l/ݙ�   3����   ���   ���   ��=���   ��=���   � >���   �>���   �>���   �>���   �������������8��������SV�t$Wjj��h � @���7����؄�tn���   P���'���؄�tZ���   Q���%���؄�tF���    ��tj�w%�����   Rj���W%���j �^%���؄�t݇�   �����$��&���؋��,P����u	_^��[� _^��[� �����̃�SV�t$W���D$P�L$Q�   h � @�Ή\$�D$    �]^����u_^3�[��� 9\$u�   R�������؄�t���   P������؄��D$    t+�L$Q������؄�t�D$��t���   RP���o���؃|$ ~��t���   W�������؋���Q����u2�_^��[��� ��������̋D$h�AP�A,�����   � �����̸m�����������V�t$��th n���������t��^�3�^���������������̸ n�����������V�t$��th�n��������t��^�3�^���������������̸�n�����������V�t$��th�o���{�����t��^�3�^���������������̸�o�����������V�t$��th�p���;�����t��^�3�^���������������̸�p�����������V�t$��th�q���������t��^�3�^���������������̸�q�����������V�t$��th�r��������t��^�3�^���������������̸�r�����������VW�|$W���B �G�F�O�N�W�V�G�F�O�N�W�O$�V�G Q�N$�F ��'���W(R�N(��'���G,�F,_��^� ���V�t$��thps��������t��^�3�^���������������̸ps�����������j�hH�d�    PQSUV�  3�P�D$d�    �L$� ��3��ωt$� ����;�~|�^V���� ��f= t"V��� ��f=
 tV��� ���L$P��(���?j�L$��(��j
�L$��(���E�;�}"S���x ��f= tS���j ��f=
 u��������;�|��L$Q�L$(��$���L$���D$�����#���ËL$d�    Y^][�����������������U������4S�]VW���i����t�   _^[��]Ë��������u���T$���T$�$踝����؍{��躜����t��诛�����D$t�D$ �s0��藜����t��茛�����D$t�D$ ��H���t�����t���i������D$t�D$ �|$ t#��蝙���%�$����4����Au��������|$ t#���s����%�$����4����Au��藙���|$ ��  ���E����%�$����4����Au���i����|$ ��  W���&�����V�\$���������T$ ��4�D$������Az[���������P  W�D$,SP�D������P�V�H�N�P�V�H�N�P�΃��V�����M�d���   _^[��]���������u	�����Y  ������Az|��������AusW�؍D$,SP�Κ�����P�V�H�N�P�V�H�N�P���ΉV�r������  ���\$ ����A��  �MSQ��d���M�d���   _^[��]�����������A�Z  S�D$,VP�N������P�W�H�O�P�W�H�O�P���ωW������t�W�D$,SP�������P�V�H�N�P�V�H�N�P���ΉV趗���M�nc���   _^[��]À|$ �  �|$ ��   V�D$,WP谙�����P�S�H�K�P�S�H�K�P���ˉS�T�����W��t��������4����A�e  ����諌�����$���V�D$,WP�H������P�S�H�K�P�S�H�K�P�˃��S�����M�b���   _^[��]�W���P������ɖ��V�D$,WP�������P�S�H�K�P�S�H�K�P���ˉS葖���M�Ib���   _^[��]À|$ t[V���������g���S�D$,VP苘�����P�W�H�O�P�W�H�O�P�σ��W�/����M��a���   _^[��]�����T$���\$���$�b�������T$����\$�$�I�������\$�����T$�$�0����M�a��_^�   [��]�������������3��y����������5���������̋A������������̃yu
�D$���   � ������������̃yu���   �3�øXt�����������j�hx�d�    P��V�  3�P�D$d�    ��t$�q����D$P�Xt�D$(    �B�������N�P�V�H�N�P�V� 0�F�0�N�0�V �0ݖ�   �F$ݞ�   �F(   �ƋL$d�    Y^�� ����軸������������SV�t$Wj j��h � @���7����؄�t.݇�   �����$�>���؄�t݇�   �����$�%���؋��lE����u	_^��[� _^��[� �����̃�SVW�|$��D$P�L$Qh � @���D$   �D$    �S���|$��t2��(��t$���   R���	���؄�t���   V���	���؋��rG����u_^��[��� _^��[��� �����̋D$h\BP��!�����   � ������݁�   ��$�5�$��������������U����j�h��d�    P��(  SVW�  3�P��$8  d�    ��t$ ��]���$���f�����  ���    ��$�   �S��$�   Ǆ$D      �d�����D$�  �t$ S���}< �������D$��   �~W�D$@P�������N(Q�T$XR������P�D$(P������L$$Q�L$@葢����;������uV��@��V�T$XR��谌��P�D$pP�������L$$�P�T$(�H�L$,�P�T$0�H�L$4�P�D$$P�L$@�T$<�,�����;�    �ٍ�$�   �����z:��$������4��������z�L$ ݁�   ��������z
ݙ�   ����؍�$�   Ǆ$@  ����������D$��$8  d�    Y_^[��]� ����$8  d�    Y_^[��]� ���̋D$���   � ��̋��   ����������j�h�d�    PQV�  3�P�D$d�    ��t$�6 ��B��=�F��=�N� >�V�>�F�>�N�>jj1�N$�D$    �V�F    �N��h�B�N(�D$�����F,    �ƋL$d�    Y^�����j�h�d�    PQV�  3�P�D$d�    ��t$��B�N(�D$   ����N$�D$ ������D$�����&6 �L$d�    Y^�������̃��x�����u�D$��thCP�����3�� �   � �V��W�N$�t���|$Ph,CW��������V�����h�&W�����_^� ���VW�|$j ��j���������tV�FP���������tD�N Q���������t2�V$R���W������t �F(P���E������t�N,Q�������_^� ����������̃�SVW���_$������t$�D$P�L$Q���D$    �D$    ����|$��u`��t^�WR��� ������tL�G P���������t:S����������t+�O(Q����������t��,W������_^��[��� 3�_^[��� ���̸    ����������̋T$3�9D$����P�D$RPQjjj j�[����� ��� ���������������̸@u�����������j�h8�d�    PQV�  3�P�D$d�    ��t$�LC���   �D$    �/�����D$�����`����L$d�    Y^������������������V�������D$t	V��������^� ��j�hv�d�    P��V�  3�P�D$d�    ��t$豮�����   �D$$    �LC�x���D$P�@u�D$(�������N�P�V�H�N�P�V� 0�F�0�N�0�V �0�F$�F(   �ƋL$d�    Y^�� �̋L$h�C�����   � ����������VW�|$��t5hHk���������t%�t$��thHk���������tW������_�^�_2�^�������������j�h��d�    P��V�  3�P�D$d�    ��t$葭�����   �D$$    �DA�(����D$P�Hk������N�P�V�H�N�P�V� 0�F�0�N�0�V �0�ΉF$�F(   ������ƋL$d�    Y^�� ����������������V���DA�2����D$t	V��������^� ������������VW�|$��t5h0l��������t%�t$��th0l��������tW���f���_�^�_2�^�������������j�hدd�    P��V�  3�P�D$d�    ��t$�Q������   �D$$    ��A�x����D$P�0l�y�����N�P�V�H�N�P�V� 0�F�0�N�0�V �0�ΉF$�F(   �b����ƋL$d�    Y^�� ����������������V����A�����D$t	V�������^� ������������V�t$��thm���k�����t��^�3�^����������������SU�l$VWU����/ �E�C�M�K�u�{�    ���   �R���   �������   ���   V������V�W�V�W�V�F�W�@�O�A���   ���   ���   ���   ���   ���   ���   ���   ���   ���   _݅�   ^ݛ�   ���   ���   ]��[� ����VW�|$��t5h�n���j�����t%�t$��th�n���R�����tW�������_�^�_2�^�������������VW�|$��tMh�o��������t=�t$��t5h�o��������t%W������݇�   ݞ�   �݇�   _ݞ�   ^�_2�^�����VW�|$��t5h�p��������t%�t$��th�p��������tW���F���_�^�_2�^�������������VW�|$��t5h�q���j�����t%�t$��th�q���R�����tW�������_�^�_2�^�������������j�h�d�    PQ�  3�P�D$d�    j0������D$���D$    t���n����L$d�    Y���3��L$d�    Y���������������j�h;�d�    PQVW�  3�P�D$d�    ��j0������D$���D$    t����������3����D$����tW��������ƋL$d�    Y_^���������������VW�|$��t5h�r���*�����t%�t$��th�r��������tW���v���_�^�_2�^�������������VW�|$W���������   ���   ݇�   ݞ�   ��݇�   _ݞ�   ^� �������VW�|$��t5hps��������t%�t$��thps��������tW������_�^�_2�^�������������U��M�T����u�D$��thDP������3�]� S���   V3���W~!3��d$ ���   �蓈����t!����;�|�m�E���w+_^[�   ]� �D$��t.h�CP�����_^[3�]� �D$��tUh�CP�{����_^[3�]� ���������������U����j�hk�d�    P���  SVW�  3�P��$�  d�    ����M���$�|�����D$J��
  �s�    ��$�   �t$`󥋃�   3�����$   ��
  �EP��$�   �V�����{
  h��jj��$p  Q�D$Z����h��jj��$H  R����h��jj��$(  P����h��jj��$   Q�n���h��jj��$�  R�X���h��jj��$�  P�B���h��jj��$p  Q�,���h��jj��$�  R����݃�   �\$L�D$K ���0c ܋�   ���$����a ܋�   ����$t  �$�����D$L��$��$�T$T��b ܋�   ���$�D$\�a ܋�   ����$�  �$�φ���D$L�b ܋�   ���$�D$T�qa ܋�   ����$�  �$虆���t$T�|$J �T  ���   ƍ�4�  P���|��݄4�  ���\$��$D  ��$Q�L$t�N����L$T��d  �P��d  �Q�P�Q�P�Q�P�Q�@Q�A��$8  Q�M�	����L$T��<  �P��@  �P��<  �Q�P�Q�P�Q�P�Q��4�  Q��4�  R����̉�P�Q�P�Q�P�Q�P�@�Q�A��$�   �N����u�D$J�ܤ4�  ����4��������{݄4�  ܤ4�  ��������Au	����D$K�D$T������`�D$T�����3���$L  �L$L�t$T3����t$T�|$J ��  ݄<l  �L$`���\$��$D  ݄<t  �$R�L�����4  �P��4  �Q�P�Q�P�Q�P�Q�@Q�A��$8  Q�M������4�  �H��4�  �P��4�  �V�H�N�P�V�H�N��<�  Q��<�  R����̉�P�Q�P�Q�P�Q�P�@�Q�A��$�   �$M����u�D$J��$�   Q��������T$L�݄<d  ܤ<�  ����4��������{݄<l  ܤ<�  ��������Au�D$K������Au	���D$J �3݃�   �xD������z���݃�   ��4������Au�D$K�D$T�D$L������H�D$T�W����|$J ��  �|$K ��  ��$�   P�L$hQ��$�  �z���L$d������$�   R��$�  P��$  �sz����$�  ������$�  Q�T$hR��$  P�݁������$  �^���\$L��$  �����$�   Q��$�  R��$,  �z����$�  �f����$�  P�L$hQ��$$  R�|�������$  ��~���\$T��$  �-���D$L�D$T������A����   ��������A��   �D$d�ًL$h�؋T$l��$�   �D$p��$�   �L$t��$�   ��$  ��$�   �T$x��$�   ��$   ��$�   ��$(  ��$�   ��$$  ��$�   ��$,  ��$�   ��$�   ��$0  ��$  ��$�   P��$  ��$�   �%y����$����z��$�   �~����$�   Q��$�   R��$<  P�   ��������A�w  �D$d�L$h�T$l��$�   �D$p��$�   �L$t��$�   �T$x��$�   ��$  ��$�   ��$  ��$�   ��$  ��$�   ��$  ��$�   ��$  ��$�   ��$  ��$�   ��$�   ��$�   P��$�   ��$�   Q��$<  R������$�   �P��$�   �H��$�   �P��$�   �H��$�   �P����$�   ��$�   �}����$�   ��H����$�   P��$8  Q��$,  �w����$�   R��$8  �w���\$L��$�   P��$8  �w���D$L��l �T$T��������Au���H+�\$T��D$J �O  ��݄$T  ܄$L  ܄$\  �5���\$|�pD�T$L��ܛ�   �����   ���   �؃�0�����tg���   �@8�@0�Fl ��������Au
���H+��݃�   ������z�����pD�*��ܳ�   ������z�������������z�����D$L�M�L$TQ���\$P�% �D$|�|$`ݓ�   ���D$d�    ݛ�   ��$�   ����\$�$���   ����~�����   ݃�   �� �Z ܋�   ���$݃�   �dY ܋�   �����$�~�����   �D$L��0�oZ ܋�   ���$�D$T�*Y ܋�   �����$�W~�����    tY���   ��$<  �SR��$D  S���ĉ��$d  �P��$h  �H��$l  �P��$p  �H��$�   �P��F���e݃�   ���   ��$�T$|��Y ܋�   ���$݄$�   �X ܋�   �����$�}����EP���"$ �|$`�    ��$�   󥍌$�   Ǆ$   �����i����D$J��$�  d�    Y_^[��]� ����$�  d�    Y_^[��]� ̋D$����|;��   }����   �����T$�L$�$�����L$���P�Q�P�@�Q�A����� �����������V��FW�|$P����I �NQ����I �VR����I ���   P���	J ���   �����P���J h�7���*J ���   Q���+J _^� ������V��F��t!��t�D$��th�EP�����3�^� W�|$W�������u��thHEW�� ����_3�^� ���   ��t��tPhEW�� ����_3�^� ���   � �X����D{2����   ���   ����\$�F�$h�DW�} ����_3�^� ���   �@ �X0����D{/��tf���   �F ���\$�F0�$hxDW�; ����_3�^� ���   �@�X8����D{/��t$���   �F���\$�F8�$h8DW�������_3�^� _�   ^� �����U������0SUVW��   3�9��   ��  ���   �sz������  ���   �� �]z������  �k�^���F����uS���������9��   ~9��   �   |���   ���   P�L$�p���L$�et�������   �؃��D$0�L$8�\$�   �D$(�$Q���&B�����H�K�P�S�H�K�P�S�@�ˉC�B���L$��r��3����L$Q���   ��o������P|���   ���T$�$��y����~���  ���   �R �J ����At�R(����D��   ��E�   �����z�B(����4����Az�Z(��   Q�؍L$�o���L$�-r���\$�L$�Pr���D$S�VXR���\$���D$8�$�J���D$ 3����T$ ��d$ �D$ ���   ���A�����D$(�����������\$�������$�y������P|���   ���T$�$��x����   ���\$�D$ �� �$��x�������t�   �F   ���   ��Y����D{
��   �Y���   �A �Y0����D{�A �   �Y0���   �@�����$�Ef�����������   u=�@8��0�$�   �"f������u���   �@(�@��$�X8���   �@8�X�S�@8��0�$��e������u���   �@�X8�+���   �A8�Y����D{�A�A8��$�Q���   �Y8�   ���    t&���   ��@�.w����u�   ���   ���    uI���   �A�YH����Dz�A0�A��$�Y@����D{ �A�   �YH���   �F0�F��$�^@���B����uS�   �G�������_^][��]Ë�_^][��]�_��^][��]�������U����j�h��d�    P��h  SVW�  3�P��$x  d�    �ى\$��M���$��������D$�q  �s�    ��$L  󥋛�   3�����$�  �  �EP��$P  �E������  h��Sj��$�  Q�D$&�!���h��Sj��$�   R����h��Sj��$  P�����h��Sj�L$@Q�����D$ 3ۀ|$ ��  �T$���   ƍ�4�   P���k��݄4  ���\$�L$,��$Q�L$,���=������  �P���  �Q�P�Q�P�Q�P�Q�@Q�A�L$ Q�M��������   �H���   �P���   �H���   �P���   �H���   �L4<Q�T48R����̉�P�Q�P�Q�P�Q�P�@�Q�A��$l  �>����u�D$��d44����4��������{݄4  �d4<��������Au	����D$������x������|$ tK�M�\$Q���; �|$ �    ��$L  �{�t$3�����   �T44R��j������P|���_�����$L  Ǆ$�  �����X����D$��$x  d�    Y_^[��]� ����$x  d�    Y_^[��]� ���   |���   � �` ������������V��F��t!��t�D$��thXFP������3�^� W�|$W�y�����u��thFW������_3�^� ���   ��t��tVh�EW�a�����_3�^� _�   ^� ����������������V�񃾘   |%���   �؍AP�D$P�������l���~u��^���������[��������������j�h˰d�    PQ�  3�P�D$d�    h�   �������D$���D$    t���[����L$d�    Y���3��L$d�    Y������������j�h��d�    PQVW�  3�P�D$d�    ��h�   �������D$���D$    t����������3����D$����t W���]���݇�   ݞ�   ݇�   ݞ�   �ƋL$d�    Y_^����VW�|$��tMhXt��������t=�t$��t5hXt��������t%W�������݇�   ݞ�   �݇�   _ݞ�   ^�_2�^�����V���B�����D$t	V���������^� ������������U������4SV��~Wt$�E����  h<IP�6�����3�_^[��]� �}W�������u!���R  h IW������3�_^[��]� ���   ��t"���&  Ph�HW�������3�_^[��]� ݆�   ���$��^��������  ��ܞ�   ������  �H+ܞ�   ������  ݆�   ���$�^�������c  ��ܖ�   �����N  ���   �A������Dz/�A������Dz#�����o  hpHW�%�����3�_^[��]� �A ������Dz/�A(������Dz#�����4  h HW�������3�_^[��]� �A0�Y0������Dz-�A8������Dz#����  h�GW������3�_^[��]� �؋��@�@�\ �\$0���   �@(�@ �\ �\$ ���   �@8�@0�q\ �T$(���D$0���������H+z���D$ ������Az��������A{��T$ ��������z��������{����\$(�������݆�   ����݆�   ��4��;������z:��t)���\$݆�   �$h�GW�������3�_^[��]� ��3�_^[��]� S�؍L$4�od�����g����ܦ�   ��݆�   ��4��;������z-��t����\$݆�   �$h@GW�T�����3�_^[��]� ���D$ �\$(����z��tph�FW�&�����3�_^[��]� �   _^[��]� �؅�tC݆�   ���$h�FW�������3�_^[��]� ��t݆�   ���$h�FW�������_^3�[��]� ������U����j�h+�d�    P��   SVW�  3�P��$�   d�    ���|$(݇�   ���$�D$/ �[�������f  ��4ܟ�   �����O  ݇�   ���$�O[�������3  ��ܟ�   �����   �H+ܟ�   �����	  �w���Pl������  �O(�@l������  �O@�0l������  �_X���l������  ���_i���%�$����4����A��  ���   ��  ���   �GV�D$@P���\$��$�   �G�$Q���n4������c���L$<��h���%�$����4����A{�L$<� i�����7  S�L$@��c������4����A�  �T$<R�D$XSP�k�����L$T�h���%�$����4����A{�L$T��h������   �]�T$@�D$D�    ���L$<�K�L$H�S�T$L�C �D$P�K$�L$T�K0�L$`�S(�T$X�S4�T$d�C,�D$\�C8�D$h�K<�S@�ˉCD�4���t$(��݆�   �L$<�\$���$�n������̉�P�Q�P�@�Q�A��Ǆ$�       ��� �L$,Ǆ$�   �����2���݆�   ݛ�   �D$'�D$'��$�   d�    Y_^[��]� �����U������8VW�}W��������   ~���   �؃�����T$�L$@�$��m����L$ �P�T$$�H�L$(�P���D$8��P�T$H��d��j ����B ���   ~���   �� �����T$�L$@�$�sm����L$ �P�T$$�H�L$(�P���D$8��P�T$H�yd��j���B ���   ~���   ��0�����T$�L$@�$�m����L$ �P�T$$�H�L$(�P���D$8��P�T$H�d��j���DB ���    ~���   �����T$�L$@�$�l����L$ �P�T$$�H�L$(�P���D$8��P�T$H��c��j����A ݆�   ݟ�   ݆�   ݟ�   _^��]� �����������W���t�D$��th�IP������3�_� V�t$V�������u��th�IV�������^3�_� ���   ��t��tWhpIV������^3�_� ^�   _� ���̃��    ���   u�@� ��@�`�����U����j�hX�d�    P��   SVW�  3�P��$�   d�    ���L$T�Ӥ���u���]Ǆ$�       tC��E�\$T�L$T�C�\$\�C�\$d� �\$l�@�\$t�@�\$|��i����u�L$T�-���3����   ��u4���   � V�@���\$�D$P�O�$P��/��P�L$\�ë���   ���uV��W�L$\誫���   ���t+�D$T�E��D$\�[�D$d�[�D$l��D$t�X�D$|�X�L$TǄ$�   ����耤���Ƌ�$�   d�    Y_^[��]� ������U����j�h��d�    P���   SVW�  3�P��$�   d�    �ًuV�S���݃�   ݞ�   �s�    �|$��݃�   ��$�   �$P�(J����$�   �$Q�L$\Ǆ$      ��]������]��P�L$�\]���L$�3/���M�T$R��3 �L$Ǆ$   ����蒣����$�   d�    Y_^[��]� ����������W���t�D$��th�JP�$�����3�_� V�t$V�������u��thhJV�������^3�_� ���   ��}��tWh0JV�������^3�_� ^�   _� ����V���(����D$t	V���������^� ��j�h��d�    PQ�  3�P�D$d�    h�   ��������D$���D$    t��������L$d�    Y���3��L$d�    Y������������j�h�d�    PQVW�  3�P�D$d�    ��h�   �Q������D$���D$    t���W������3����D$����tW�������Ǹ   W���   �����ƋL$d�    Y_^����������VW�|$��tGh@u���ʷ����t7�t$��t/h@u��買����tW��覃���Ǹ   W���   �D���_�^�_2�^����������̃�V�t$��t4�D$P�@u�Ŵ��P���M�������th@u���K�����t��^���3�^������������j�h�d�    PSVW�  3�P�D$d�    �|$ ����   W�{����\$(���ۋ�t_f�; tY��u6h�   ��������D$ ���t$t	��������3�P���D$�������.���S���   ������L$d�    Y_^[��Å�t��Pj���ҋL$d�    Y_^[���������������̃�V���t=�D$P�@u觳��P���/�������t h@u���-�����t���   �~���^���3�^�����j�hK�d�    PQ�  3�P�D$d�    h�   ��������D$���D$    t�������L$d�    Y���3��L$d�    Y������������j�h{�d�    PQVW�  3�P�D$d�    ��h�   �������D$���D$    t���������3����D$����tW���}����ƋL$d�    Y_^������������j�h��d�    PQ�  3�P�D$d�    h�   �������D$���D$    t���k����L$d�    Y���3��L$d�    Y������������j�h۲d�    PQVW�  3�P�D$d�    ��h�   �������D$���D$    t����������3����D$����tW���-����ƋL$d�    Y_^������������VW�|$��t5h n��������t%�t$��th n��������tW������_�^�_2�^�������������SU�鋅�   3�;�VWt���   ��QSP�' �����   S�Ή��   �����3��F�FS�FU�F�a������]�}�    �hY�_^���   ���   ƅ�   ][�����j�h/�d�    PQSVW�  3�P�D$d�    ���|$��J�D$   �C������   �D$�#������   3�9^�D$�lIt�F;�tSP���xI�^�^�^�O�\$�Ŝ�����D$�����v �L$d�    Y_^[�����̃�(SV��L$4�A���2ۃ�wl�AP�L$Q���H����L$��^����tO�D$���\$�T$(�D$�N�$R�,'����L$8��P�Q�P�Q�P�Q�P�Q�@^�A�[��(� ����D$8�����P����H����P����H����P^��[��(� ���������j�hX�d�    P��SUVW�  3�P�D$$d�    ��������|$43���Ɔ�    �D$ �D$�֪����|4���J>  =$��|&�D$P�L$$Qh � @���D$@������u'3���  �T$R�D$$P���D$< �'����؄���  �|$ t2��  �L$Q���#����؄���  �T$R�����F���D$P��������؄��z  �L$�V�NR���!����؄��^  ���   U��������؄��F  ���   P�������؄��.  �L$Q���D$    �����؄��  �|$ ���   ��P�ψ��   �m����؄���   ���   Q��������؄���   �F����   ;�w.�$�n���   }%����    ����   u9M|�MƆ�    �|$4 ��   ���   R��������؄�to�D$��~g��|b���   P���-����؄�tN�|$|G�L$�����D$P���D$0    �����؄ۍL$t�����PV�]������L$�D$,���������|$4 t��������u2��ËL$$d�    Y_^][��� mm&m1m1m��������U����j�h��d�    P��   SVW�  3�P��$�   d�    ��L$T�C����]�ۋ}Ǆ$�       tC��E�\$T�L$T�G�\$\�G�\$d� �\$l�@�\$t�@�\$|�Z]����u�L$T蝘��3ۋ��   ���S  P�L$ ����L$,Ƅ$�   ��P�����    t4���   � ���T$<�N�@�D$L�T$D�\$�$P�#��P�L$ �=���~W�L$ �w=����   �T$,�A���T$D�T$L�\$���$R��"��P�L$ �D=�����   �@ �� �T$,���@�D$L�T$D���\$�$P�"��P�L$ �=�����   �A���T$D�T$L�\$���D$<�$R�f"��P�L$ ��<��S�D$pP�L$\Q�L$(�����|$( ��Ƅ$�    �D$�$t"�D$ ��t3�VP�L$$��$�t$ �t$(�t$$�}��t+�D$T�E��D$\�_�D$d�_�D$l��D$t�X�D$|�X�L$TǄ$�   ���������Ë�$�   d�    Y_^[��]� ������������U����j�hȳd�    P��hSVW�  3�P�D$xd�    �����   ����   P�L$ �ɑ��3���$�   �_���   �D0ƃ��\$�L$<� �$Q���)!��P�L$ �;������P|ʋU�u�ERVP�L$(�E ��t�   �|$( Ǆ$�   �����D$�$t5�D$ ��t-j P�L$$��$��u��t�}���Z����u	���ܕ��3�3������L$xd�    Y_^[��]� ��������������U����j�h�d�    P��   SVW�  3�P��$�   d�    ��L$T�Ô���]�ۋ}Ǆ$�       tC��E�\$T�L$T�G�\$\�G�\$d� �\$l�@�\$t�@�\$|��Y����u�L$T����3ۋ��   ���]  P�L$ �B����L$,Ƅ$�   �AM�����    t4���   � ���T$<�N�@�D$L�T$D�\$�$P���P�L$ �:���~W�L$ ��9�����   �@���T$,���@�L$L�T$D�\$�$Q���J��P�L$ ��9�����   �@ �� �T$,���@�T$L�T$D���\$�$R���P�L$ �9�����   �F0��0�T$,���F�D$L�T$D���\$�$P����P�L$ �R9��S�L$pQ�T$\R�L$(�~����|$( ��Ƅ$�    �D$�$t"�D$ ��t3�VP�L$$��$�t$ �t$(�t$$�}��t+�D$T�E��D$\�_�D$d�_�D$l��D$t�X�D$|�X�L$TǄ$�   �����\����Ë�$�   d�    Y_^[��]� ��U����j�h8�d�    P��hSVW�  3�P�D$xd�    �����   ����   P�L$ �I���3���$�   �_���   �D0ƃ��\$�L$<� �$Q�����P�L$ �8������@|ʋU�u�ERVP�L$(�B ��t�   �|$( Ǆ$�   �����D$�$t5�D$ ��t-j P�L$$��$��u��t�}���W����u	���\���3�3������L$xd�    Y_^[��]� ��������������U����j�hv�d�    P���   SVW�  3�P��$�   d�    �L$�L$�A����u���}�]Ǆ$�       t@��L$�\$�G�\$�G�\$$��\$,�C�\$4�C�\$<�XV����u�L$蛑��3��L$D�� �L$�D$DPƄ$�   ������t#3Ʌ���j �T$QR�L$P�J ��t�   ���t(�D$��D$�_�D$$�_�D$,��D$4�[�D$<�[�L$DƄ$�    �f� �L$Ǆ$�   ���������Ƌ�$�   d�    Y_^[��]� ��������j�h��d�    P��   SVW�  3�P��$�   d�    ��L$��� �D$P��Ǆ$�       ��������$�   t%��$�   ��$�   QVR�L$�-I ��t&�   ���t��$�   ��� U����u	���E���3����L$��Ǆ$�   �����z� �Ë�$�   d�    Y_^[�Ĥ   � ������������̃�V�t$W3����ΉD$�D$�$�����|7���2  =$��|)�D$P�L$Qh � @���D$ �&����u_3�^��� �D$ SV���������Ä�t$���   R�������؄�t���   W��������؀|$ t��������u2���[_^��� ������������̃�UV�t$W���D$P�L$Q3�h � @�Ήl$�l$�������   �|$St2��   �T$R�D$$Ph � @�Ήl$,�l$$�O���؄�t;�|$ t2��V����������Ë��:����u2����t���   Q��������9l$~(��t$���   R�������؄�t���   W�������؋�������u[_^��]��� ��[_^]��� _^��]��� ���������������U����j�h�d�    P��   SVW�  3�P��$�   d�    ��L$T�C����]�ۋ}Ǆ$�       tC�E� �L$T�\$T�@�\$\�@�\$d��\$l�G�\$t�G�\$|�ZR����u�L$T蝍��3ۋ��   ����   P�L$0������   �@���\$�~� �D$L�$P��Ƅ$�   �&��P�L$0�2�����   �F���\$�L$L�F�$Q������P�L$0�p2��S�T$pR�D$\P�L$8蜀���|$8 ��Ƅ$�    �D$,�$t"�D$0��t3�VP�L$4��$�t$0�t$8�t$4�}��t+�E�D$T��D$\�X�D$d�X�D$l��D$t�_�D$|�_�L$TǄ$�   �����z����Ë�$�   d�    Y_^[��]� U����j�h�d�    P��lVW�  3�P�D$xd�    �񋆘   ����   P�L$ �j������   �@���\$�~� �D$<�$P��Ǆ$�       ����P�L$ �A1�����   �F���\$�L$<�F�$Q�����P�L$ �1���U�u�ERVP�L$(�; ��t�   �|$( Ǆ$�   �����D$�$t5�D$ ��t-j P�L$$��$��u��t�}���P����u	���Z���3�3������L$xd�    Y_^��]� �������������U��}t�D$��thLNP�������3�]� SV���   W���������3���~�I V������f=  w<��;�|��}���o�����tf�8 u�D$��t9hNP�r�����_^[3�]� �t$V���:�����u��th�MV�G�����_^[3�]� ���   ��t��tUh�MV�!�����_^[3�]� _^[�   ]� ��������̃�V�t$W3����ΉD$�D$�d�����|7����,  =$��|)�D$P�L$Qh � @���D$ �f	����u_3�^��� �D$ SV����������À|$ t���G�����u2���[_^��� �����j�hH�d�    P��(VW�  3�P�D$4d�    �񋆘   ����   P�L$谄�����   �@���\$�N� �D$,�$P�D$P    ���P�L$�.���L$L�t$H�T$DQVR�L$�8 ��t�   �|$ �D$<�����D$�$t7�D$��t/j P�L$��$� �t$H��t�|$D���M����u	���ψ��3�3������L$4d�    Y_^��4� ��U����j�h��d�    P��   SVW�  3�P��$�   d�    ���L$T�Ç���u3�9]��$�   tD��E�\$T�L$T�F�\$\�F�\$d� �\$l�@�\$t�@�\$|��L����u�L$T�!����]���   ����   S�L$0�F�����Ƅ$�   ~D3����    ���   �0��@���\$�D$L�O�$P���P�L$0�-������uɋu3�9M�T$T��QR�L$4�?�����t�E   �|$8 Ƅ$�    �D$,�$t"�D$0��t3�WP�L$4��$�|$0�|$8�|$4�}��t+�D$T�E��D$\�^�D$d�^�D$l��D$t�X�D$|�X�L$TǄ$�   ���������ǋ�$�   d�    Y_^[��]� �����������U����j�h��d�    P��hSVW�  3�P�D$xd�    �����   ����   S�L$ ����3�;މ�$�   ~7���   �0��@���\$�D$<�O�$P�G��P�L$ �+������uɋM�u�UQVR�L$(�5 ��t�   �|$( Ǆ$�   �����D$�$t5�D$ ��t-j P�L$$��$��u��t�}���J����u	�������3�3������L$xd�    Y_^[��]� ������������j�h�d�    PQVW�  3�P�D$d�    ��t$��� �N�D$    ��J�������   �D$�������   ���D$�Z���3��G�G�G�G���ݞ�   �D$�F   ǆ�   �����W����ƋL$d�    Y_^������V�������D$t	V��������^� ��j�h@�d�    P��SUVW�  3�P�D$,d�    ��t$<�������������D$<��tjjh � @�.l����u3��2  3�Wj�Y����؄��  �3��EP�������؄���  �EP���k����؄���  �EP���&����؄���  ���   Q�L$ ����E3�8��   �   ���;��|$4�T$ws�$���9L$$uj�L$�ԯ���D$ �@���\$�H@�@ � ��$�$��F���79L$$u	�L$蟯���|$$|!�L$ �Q �A ��@��P�Q�P�Q�@�A�|$�L$Q���w����؄���   ���ƒ�������   V腧��������   R�������؄���   �D$P���L����؄���   ���   Q���4����؄���   ݅�   �����$�����؄�tx�|$< u�L$�D$4��������   ���   R��������؄�tG���   P�������؄�t2���d���P�L$������L$Q���D$8�Y����L$���D$4 �����L$�D$4�����(���|$< t���j�����u2��ËL$,d�    Y_^][��$� �I =�=���r�r�����U����j�hv�d�    P��h  SVW�  3�P��$x  d�    �ى\$(��M���$��������  ���    ��$�   �EP��$�   Ǆ$�      �R�����D$&�1  �|$(���   V�L$8�t$0�>|����$�   Ƅ$�  ��9���L$D��9���L$T��9����$�   �9�����D$' �D$0    �{  3���I �|$& ��  ���   �0�ݔ$�   ���@�L$|ݔ$�   �\$�$Q��������T$T�H�L$X�P�T$\�H�L$`�P�T$d�@�L$TQ�M�T$pR�D$p��������$�   �P��$�   �H��$�   �P��$�   �H��$�   �P��$�   �L$LQ�T$HR����̉�P�Q�P�Q�P�Q�P�@�Q�A��$�   �P����u�D$&݄$�   �D$D������4��������u���\$D����D$'݄$�   �D$L������������Az�\$L����D$'�L$DQ�L$8�X���D$0����;D$,�D$0������|$& �  �UR���F� �|$' �    ��$�   ���|$(t�D$4P���   �z����   �����Dz�Y����D��   ���Q�L$p��7���L$l�E<������   �D$t���\$��$�   �D$|�$Q���
�����H�K�P�S�H�K�P�S�@�ˉC�
���L$l��:���D$,��~+�   �X����$    �L$lQ���   ��7������u���   ���T$�$�A���|$@ Ƅ$�   �D$4lIt#�D$8��tj P�L$<�xI3��D$8�D$@�D$<��$�   Ǆ$�  �����^~���D$&��$x  d�    Y_^[��]� ����$x  d�    Y_^[��]� ������j�h��d�    PQSVW�  3�P�D$d�    �ى\$�1����DK�C   �C   �{�    �hY󥍳�   hB���D$     �����3��F�FP�FS�F�������   ���   �   ��;�}O9~~�~�N��PWQ���҅��Ft$�N;�}��+���R���j Q� ���~��F    �F    9~|�~�F��t�v��~��Vj P�v ���ËL$d�    Y_^[�����������������V���DK�����D$t	V���������^� ������������SV�t$W����� ������Ä�tj jh � @���&d����u_^3�[� V���������D$��t���p�����u�D$�D$_^[� �������������j�hضd�    PQSVW�  3�P�D$d�    ���|$�a������   �   hD���D$     ��K�_�G   �"���3��F�FP�FW�F�������   ���   ��;�}O9^~�^�N��PSQ���҅��Ft$�N;�}��+���R���j Q�� ���^��F    �F    9^|�^�F��t�v��~��Vj P� ���ǋL$d�    Y_^[����V����K������D$t	V�E�������^� ������������j�h�d�    PQSVW�  3�P�D$d�    ��t$�!�����ݞ�   ���   ��hB��ݞ�   �D$     �4L�F   �F   �����3��G�GP�GV�G�n������   ���   �   ��;�}O9_~�_�O��PSQ���҅��Gt$�O;�}��+���R���j Q� ���_��G    �G    9_|�_�G��t���~��Wj P�e ���ƋL$d�    Y_^[����������������V���4L�����D$t	V���������^� ������������V�t$W���������������D$tj jh � @���a����u_3�^� SV���������Ä�t.݇�   �����$�����؄�t݇�   �����$������؀|$ t���*�����u2���[_^� �����������j�h8�d�    PQSVW�  3�P�D$d�    ���|$�!������   hB���D$     ��L�G   �����3��F�FP�FW�F�������   Ǉ�   �����F�   ��;�}O9^~�^�N��PSQ���҅��Ft$�N;�}��+���R���j Q� ���^��F    �F    9^|�^�F��t�v��~��Vj P�u ���5��ݗ�   ݟ�   �L$d�    Y_^[��������������V����L�����D$t	V���������^� ������������V�t$Wjj��h � @���(_������   Sj jh � @���_���؄�tbV�������������e�����u2��F��tB���   P���[����؄�t.݇�   �����$�����؄�t݇�   �����$�ɾ���؋�������u	[_��^� ��[_^� _��^� ��V���$M�����D$t	V���������^� ������������V����N�b����D$t	V���������^� ������������j�hk�d�    PQ�  3�P�D$d�    h�   腿�����D$���D$    t���+����L$d�    Y���3��L$d�    Y������������j�h��d�    PQVW�  3�P�D$d�    ��h�   �������D$���D$    t���������3����D$����tW���}����ƋL$d�    Y_^������������j�h˷d�    PQ�  3�P�D$d�    h�   蕾�����D$���D$    t�������L$d�    Y���3��L$d�    Y������������j�h��d�    PQVW�  3�P�D$d�    ��h�   �!������D$���D$    t���������3����D$����tW��荪���ƋL$d�    Y_^������������j�h+�d�    PQ�  3�P�D$d�    h�   襽�����D$���D$    t���[����L$d�    Y���3��L$d�    Y������������j�h[�d�    PQVW�  3�P�D$d�    ��h�   �1������D$���D$    t����������3����D$����t W��蝩��݇�   ݞ�   ݇�   ݞ�   �ƋL$d�    Y_^����j�h��d�    PQV�  3�P�D$d�    h�   褼�������t$���D$    t.�������$M�F   �F    �ƋL$d�    Y^���3��L$d�    Y^�����������������j�h��d�    PQSV�  3�P�D$d�    ��h�   ���������t$���D$    t�������$M�F   �F    �3����D$����tS���i����ƋL$d�    Y^[��������j�h�d�    PQV�  3�P�D$d�    h�   脻�������t$3�;��D$t��������N�F   �F   �ƋL$d�    Y^������j�h�d�    PQVW�  3�P�D$d�    ��h�   ���������t$���D$    t��������N�F   �F   �3����D$����tW���i����ƋL$d�    Y_^��������j�hK�d�    PQ�  3�P�D$d�    h�   腺�����D$���D$    t���;����L$d�    Y���3��L$d�    Y������������j�h{�d�    PQVW�  3�P�D$d�    ��h�   �������D$���D$    t����������3����D$����t,W���}������   ���   ݇�   ݞ�   ݇�   ݞ�   �ƋL$d�    Y_^��������U������   S�]VWS����� �L$�(���L$@����j ���+�������$������4���������!  ����������A�  �pD�N �T$(���T$�L$X�T$�$賴��3�9��   ��   3ۍI ����|;��   }���   �������T$�L$@�$��5����L$�P�T$�H�L$ �P�D$@P�L$�T$(�%����|A���   ;�}%���   �L$É�T$�P�L$ �H�T$$�P�u�D$P���   ��G������;��   �S����]�~u%݆�   �L$(��4������z
ݞ�   �����S�N� ��_^��[��]� �k����������������VW�|$������$�������uW���=���_^� _��^� ���3ɉH��H��V�t$��th0v��蛄����t��^�3�^���������������̸0v����������̋D$�A�� ����V��~ ��Qt%�F��tj P��Q�F    �F    �F    ^�����������V��~ ��Qt%�F��tj P��Q�F    �F    �F    �D$t	V��������^� ������VW�|$��t5h0v��躃����t%�t$��th0v��袃����tW���Ƌ��_�^�_2�^�������������j�h��d�    PQVW�  3�P�D$d�    ��t$����3��N�|$��Q�F�����'���3��F �Q�~$�~(�~,�F�F�F�F�ƋL$d�    Y_^��������j�h�d�    PQSUVW�  3�P�D$d�    ���|$��Q�o���D$    �Ͱ���w 3�9^�D$ ��Qt�F;�tSP����Q�^�^�^�͈\$ 蓰�����D$ ���������L$d�    Y_^][���QS�Y(���L$}�D$��thdSP�������3�[Y� ��UVWu_��I$�����u$�D$���;  hSP�ɳ����_^]3�[Y� �y ��   �D$���  h�RP蛳����_^]3�[Y� 3���~d�i$��3ҍ}�*����At]���t��ut��t2�A$�L�;H���   �*������Dz�G�������D��   �L$������;�|���_^]�   [Y� �D$�؅�tth�RP������_^]3�[Y� �D$�؅�tRh�RP������_^]3�[Y� �D$�؅�t0hLRP農����_^]3�[Y� �D$�؅�thRP蜲����_^]3�[Y� ���������������V�t$Wjj��h � @���(R����t^�GSP��蘰���؄�t/�GP���7����؄�t�O Q��������؄�t��W���U����؋��L�����u	[_��^� ��[_^� _��^� ����������������V�q(W3���|*�A$�V����� ���<�    �@���@���@��@��@�u�;�}����A$+�� ����u�_^��������������j�h�d�    PQ�  3�P�D$d�    j0踲�����D$���D$    t�������L$d�    Y���3��L$d�    Y���������������j�hK�d�    PQVW�  3�P�D$d�    ��j0�D������D$���D$    t���������3����D$����tW���0����ƋL$d�    Y_^���������������V��������D$t	V�۳������^� ��3�V���F�����F�F�F�N�F谬���� �~ t(�F��t!�j P�B�����F    �F    �F    ^��������������SUW���O賮���G(�l$Ph�SU� ��������������$h�SU����h�SU�گ��3ۃ�9_(~U�\$V�w$t$��thKU赯�����v�� t��th�S�h�S�h�SU茯���D$����;_(|�^hKU�p�����_][� ������̃�SVW��������|$3��D$�D$�D$P�L$Q�^h � @��������������tZ�|$uFS���S����؄�t�VR���2����؄�t�F P�������؃|$|��t��V���9������2ۋ�������u_^��[��� _^��[��� �T���������̃�Q�L$����� ��Q�L$����� ��Q�L$�C���� ��Q�L$����� ��Q�L$裣��� ��Q�L$�#���� ��Q�L$����� ��Q�L$胥��� ��Q�L$�s���� ��Q�L$����� ��Q�L$����� ��Q�L$賣��� ��Q�L$�S���� ��Q�L$������ ��Q�L$������ ��Q�L$����� ��Q�L$�S���� ��Q�L$�3���� � w����������̋T$�ҋD$u���Å�u�   Ë���u��ɋ�Å�t�@+A�����������̋D$�Q ��Q$�P�Q(�I,�P�H� ��j�h��d�    PQV�  3�P�D$d�    ��t$�S� ���   �D$    � �����   �D$������   �D$� ���ƋL$d�    Y^����������������j�hԺd�    PQV�  3�P�D$d�    ��t$���   �D$   �d�����   �D$�ud�����   �D$ �ed�����D$������ �L$d�    Y^��������VW�|$j j��h � @���K����u_^� SW��2��d� ��tK���   P���Q�����t8���   Q���?�����t&���   R���-�����t���   V��������t���������u2ۊ�[_^� ��SUV3�W��D$�D$��� ���   ���   ���E  �*�����   �L$�*�����   �L$��)���|$$�D$P�L$Qh � @���������u_^]2�[��� �|$�D$$ uIW���� ��t=U��艦����t1S���-�����t%�T$R��������t�D$P��������t�D$$���m�����t��D$$_^][��� ����������̋Q2���t(�I��~!V�t$��t��~Vh@  QR�5]�����^� �����������̋Q2���t(�I��~!V�t$��t��~Vh@  QR��\�����^� �����������̋D$�L$����PQ�������� ����̋D$�L$i��   PQ������� ����̋Q2���t%�I��~V�t$��t��~VjQR�x\�����^� ��������������̋Q2���t%�I��~V�t$��t��~VjQR�(\�����^� ��������������̋D$�L$��PQ������� �������̋Q2���t%�I��~V�t$��t��~VjdQR��[�����^� ��������������̋Q2���t%�I��~V�t$��t��~VjdQR�[�����^� ��������������̋D$�L$k�dPQ�n������ ��������j�h�d�    PQ�  3�P�D$d�    �L$�L$���D$    t�F����L$d�    Y��� ����S�\$��U��~[W�|$��|QV�t$��|G;�tC�E�;�9;�5�M�;�~�;�}��P����z���E����S����WV��� ��^_][� ����VW�|$W���� ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ��   +��@   ������u�_��^� ������D$V���Tt	V�:�������^� �SUVW�|$��]h�TW�Ȧ�������>���3���~,���    �E�< �tEu�lEPW薦������;�|܋��E���_^]�[� ������������SUVW�|$�ًkh�TW�X��������Υ��3���~�C��Qht:W�6�������;�|������_^]�[� ������������U������4SVW�}�ًCh�TW�D$D���������c���3�9t$<~�K������$������;t$<|���x���_^�[��]� �������������SUW�|$�ًkh UW艥�������������~V3��C�P���K�������u�^������_]�[� ���SUW�|$hUW���<�������貤���k��~V3��C�P���ۨ������u�^���ˤ��_]�[� ��̋A�������������SUW�|$h UW���ܤ�������R����k��~V3��C�P�������ƀ   ��u�^���h���_]�[� �A�T$��A� �QSUV��W�L$耊���|$h@UW�q������������k3���~=�C���L$�L$蛊��P�L$聊��P�L$�g���Ph0UW�+�������;�|Ë��ڣ��_^]�[Y� SUW�|$hPUW������������r����k��~V3��C�P���;�������u�^��苣��_]�[� ���SUVW�|$h\UW��諣�������!����k3���~�C��Q��芪����;�|���<���_^]�[� ���SUV�t$hxUV���\��������Ң���k��~@W3����    hlUV�5����C���P��腩��h�&V���������   ��u�_���Ģ��^]�[� ������������V�t$h�UV���������V�����菢���^� ���������V�t$��th w����p����t��^�3�^����������������SV��^hW3���~$���Fd���ɍ��     t��j�Ѓ�;�|ރ~l |�Fh    �`/�N �d/�V$�h/�F(�l/�N,�F    �F    �`/�V�d/�F�h/�N�l/�N0�V�UM��_�NH^[�JM������������QUV�t$jj��h � @���A����u^3�]Y� S�E P���ߡ���؄��H  �MQ���ڟ���؄��3  �UR��赡���؄��  j V�MH�`N���؄��	  V�M0��W���؄���   j jh � @���A���؄���   W�}hW�Ή|$�i��������D$    ��   ��$    ����   j jh � @���@���؄�tt�Ed�L$�<���t�G�3�P�������؄�t/��t�G�3�P��������؄�t��t� t��BV���Њ؋��������u2ۋD$��;D$�D$�n�����������_u2����t�MQ��蟞���؋�������u2���[^]Y� ������S�\$Vj j��h � @����?����u^2�[� �FP���D$ �M�����tiW3�;~}$U3�N�S�������t����@  ;~|�;~]_|:�FP��������t+�F��~�NQP��������t�F P��������t�D$����������m����D$^[� ��������V��~ �tTt%�F��tj P��T�F    �F    �F    ^�����������V��~ �tTt%�F��tj P��T�F    �F    �F    �D$t	V�O�������^� �����̋D$9A}	�D$����� �����������VW�|$��;�t>�G��_�F    ��^� 9F}P�q���N��t�G�F��P�GPQ�)� ��_��^� ���������������V��L$��|6�F;�}/+���P�APQ�������F��F��Fh�   j P��� ��^� �����������V��~ ��Tt%�F��tj P��T�F    �F    �F    �D$t	V�/�������^� �����̋��@   �@����� �U3��@�H�H�H�H��������j�h(�d�    PQSVW�  3�P�D$d�    ���|$��U3�9_�w�\$��Ht�F;�tSP����H�^�^�^�T�L$d�    Y_^[������������j�hX�d�    PQV�  3�P�D$d�    ��t$�D$�T�H�N�P�V3ҍN��U��P�T$��H�Q�Q�Q��H�ƋL$d�    Y^��� ����̋��@   �@����� �U3��@�$�H�H�H��������j�h��d�    PQSVW�  3�P�D$d�    ���|$��U3�9_�w�\$��$t�F;�tSP����$�^�^�^�T�L$d�    Y_^[������������j�h��d�    PQV�  3�P�D$d�    ��t$�D$�T�H�N�P�V3ҍN��U��P�T$��$�Q�Q�Q��$�ƋL$d�    Y^��� ����̋��@   �@����� <V3��@%�H�H�H��������j�h�d�    PQSVW�  3�P�D$d�    ���|$�<V3�9_�w�\$�%t�F;�tSP���%�^�^�^�T�L$d�    Y_^[������������j�h�d�    PQV�  3�P�D$d�    ��t$�D$�T�H�N�P�V3ҍN�<V��P�T$�%�Q�Q�Q�%�ƋL$d�    Y^��� ����̋��@   �@����� �V3��@�$�H�H�H��������j�hH�d�    PQSVW�  3�P�D$d�    ���|$��V3�9_�w�\$��$t�F;�tSP����$�^�^�^�T�L$d�    Y_^[������������j�hx�d�    PQV�  3�P�D$d�    ��t$�D$�T�H�N�P�V3ҍN��V��P�T$��$�Q�Q�Q��$�ƋL$d�    Y^��� ����̋��@   �@����� �V3��@��H�H�H��������j�h��d�    PQSVW�  3�P�D$d�    ���|$��V3�9_�w�\$��t�F;�tSP���$��^�^�^�T�L$d�    Y_^[������������j�hؼd�    PQV�  3�P�D$d�    ��t$�D$�T�H�N�P�V3ҍN��V��P�T$���Q�Q�Q���ƋL$d�    Y^��� ����̋��@   �@����� ,W3��@�T�H�H�H��������j�h�d�    PQSVW�  3�P�D$d�    ���|$�,W3�9_�w�\$��Tt�F;�tSP����T�^�^�^�T�L$d�    Y_^[������������j�h8�d�    PQV�  3�P�D$d�    ��t$�D$�T�H�N�P�V3ҍN�,W��P�T$��T�Q�Q�Q��T�ƋL$d�    Y^��� ����̋��@   �@����� |W3��@�H�H�H�H��������j�hh�d�    PQSVW�  3�P�D$d�    ���|$�|W3�9_�w�\$��Ht�F;�tSP����H�^�^�^�T�L$d�    Y_^[������������j�h��d�    PQV�  3�P�D$d�    ��t$�D$�T�H�N�P�V3ҍN�|W��P�T$��H�Q�Q�Q��H�ƋL$d�    Y^��� ����̋��@   �@����� �W3��@�[�H�H�H��������j�hȽd�    PQSVW�  3�P�D$d�    ���|$��W3�9_�w�\$��[t�F;�tSP����[�^�^�^�T�L$d�    Y_^[������������j�h��d�    PQV�  3�P�D$d�    ��t$�D$�T�H�N�P�V3ҍN��W��P�T$��[�Q�Q�Q��[�ƋL$d�    Y^��� �����QUW�|$j j��h � @����3����u_]Y� �ESP���a����؄�t6�EV3����D$~'3���t�M�D$�P��������d;t$��|ߋ|$^��������u2ۊ�[_]Y� ���������������j�h3�d�    PQVW�  3�P�D$d�    ��t$�r_��3�j�N0�|$�X�\I��j�NH�D$�MI���F`tT�~d�~h�~l�`/�F�d/�N�h/�V�l/�F�~�~�`/�N �d/�V$�h/�F(�l/�N,�Fp�ƋL$d�    Y_^�������������j�hy�d�    PQSUVW�  3�P�D$d�    ���|$�X�_h�o`3�9u�D$    |�u;�~�Gd����t��j�Ѓ�;�|�} �D$ �E tTt�E��tj P����T3��E�E�E�OH�D$ �nH���O0�D$  �aH�����D$ ������e���L$d�    Y_^][�����������������j�h��d�    P��SUVW�  3�P�D$(d�    �ًkh3�3�3�;�t$�D$�$�L$�t$ �D$$~U�L$������L$�D$$;�t$0|;��l$ ;�t;�~��PVQ�� �L$(���Sd;�t;�Ch;�~4�����t+��t'��~h��jPRQj�5 ���u
�    �L$3���~S�t$8���Sd����t7�@PhLXV��������蓐���Kd����BV�Ћ�辐���D$�L$��;�|��t$�|$$ �D$0�����D$�$t��tj Q�L$ ��$�ƋL$(d�    Y_^][�� � ����������j�hؾd�    P��SUVW�  3�P�D$$d�    ��3��D$�[�|$�|$�|$ �t$4hYV�|$4�N������EP��蠖��h�&V�5����MQh YV�&���h�XV�������U R���m���h�&V�������}��Xt��XPh�XV������9|$ |�|$�D$P�M0��L���\$;�h�XV趏�����Gh�XV規����������;�~'�L$�R������h�&V�~���������u�3����*���9|$ |�|$�D$P�MH�sL���\$;�h�XV�@������IhpXV�0�������覎��;�~)���L$�R���q���h�&V����������u�3���貎��hdXV���������]���V�������;�uh\XV�Ǝ�������|���9|$ �D$,�����D$�[t�D$;�tWP�L$��[�L$$d�    Y_^][��� ������������SUVW�|$����}V3�9n�  �~��x%�������    �N���������@  ;�}�N��PUQ����_�n�n�n^][� �F;�}n�N��PWQ����3�;ŉF��   �V��+ʍ�����Q���UR�\� �F��;�}"������+�F�P��������@  ��u�~_^][� ~Q���;�|"��+�������N��������@  ��u�9~~�~��F�RWP�Ή~��3�;ŉFu�n�n_^][� ������������U�l$V��;�t[�ES3�;��^[��^]� 9F}P����9^t�E;ÉF~�W3����E�N�P���������@  ;^|�_[��^]� ��^]� ��V�������D$t	V���������^� ��j�h�d�    PQV�  3�P�D$d�    ��j�ō�����D$���D$    tV���:����L$d�    Y^���3��L$d�    Y^���������V�������D$t	V�k�������^� ��j�h;�d�    PQV�  3�P�D$d�    ��j�5������D$���D$    tV��������L$d�    Y^���3��L$d�    Y^���������V���X����D$t	V�ێ������^� ��j�hk�d�    PQV�  3�P�D$d�    ��j襌�����D$���D$    tV���z����L$d�    Y^���3��L$d�    Y^���������V��������D$t	V�K�������^� ��j�h��d�    PQV�  3�P�D$d�    ��j�������D$���D$    tV�������L$d�    Y^���3��L$d�    Y^���������V�������D$t	V軍������^� ��j�h˿d�    PQV�  3�P�D$d�    ��j腋�����D$���D$    tV�������L$d�    Y^���3��L$d�    Y^���������V���8����D$t	V�+�������^� ��j�h��d�    PQV�  3�P�D$d�    ��j��������D$���D$    tV���Z����L$d�    Y^���3��L$d�    Y^���������V��������D$t	V蛌������^� ��j�h+�d�    PQV�  3�P�D$d�    ��j�e������D$���D$    tV��������L$d�    Y^���3��L$d�    Y^���������V���x����D$t	V��������^� ��j�h[�d�    PQV�  3�P�D$d�    ��j�Չ�����D$���D$    tV�������L$d�    Y^���3��L$d�    Y^���������j�h��d�    PQ�  3�P�D$d�    jt�h������D$���D$    t���>����L$d�    Y���3��L$d�    Y���������������V��������D$t	V��������^� ��QSUV��W�|$�G�F�O�N�W�V�G�F�O�N�W�V�G �F �O$�N$�W(�V(�G,�OHQ�NH�F,�=���W0R�N0�=���Fp�oh�N`U�k��3�;�\$~V��$    �Gd����t>��B�Ѕ��D$t/�L$Q�N`�z����~p �L$t�D$��t�P;Q~�Fp �L$��;�|�_^][Y� ���������UW��3�9o�`Tt:V�w��xS�����O���������@  ;�}�[�O��PUQ���҉o^�o�o_]�������������V�������D$t	V諉������^� ��UW��3�9ot?V�w��x$S������I �O���������@  ;�}�[�O��PUQ���҉o^�o�o_]��������������UV��3�9n��Tt<W�~��x!S��i��   �N�裶 �����   ;�}�[�N��PUQ���҉n_�n�n^]�����������U�l$V��;�t[�ES3�;��^[��^]� 9F}P�T���9^t�E;ÉF~�W3����E�N�P��0� �����   ;^|�_[��^]� ��^]� ��SV��3�9^��Tt1W�~��x��    �F���E�����y���F�RSP���҉^_�^�^^[������S�\$V��;�tT�CW3�;��~_��^[� 9F}P�t���9~t.�C;ǉF~$��I �K��    �Q�N��i�����;~|�_��^[� ���������V���h����D$t	V蛇������^� ��V�������D$t	V�{�������^� ��VW�|$W��������F�@�N�WR�ЋO �N �F$+��@   �I ������u�_��^� �����������̋��@   �@����� $Y3��@�T�H�H�H��������j�h��d�    PQV�  3�P�D$d�    ��t$�$Y�N�D$    �B����T�L$d�    Y^��������������V��L$�FP�`����F^� ��������̋��@	   �@����� tY3��@�T�H�H�H��������j�h��d�    PQV�  3�P�D$d�    ��t$�tY�N�D$    ������T�L$d�    Y^��������������V��L$�FP������F^� ���������j�h�d�    PQVW�  3�P�D$d�    ��jt蔃�����D$���D$    t���j������3����D$����t;�t���}���W���[��W���M����ƋL$d�    Y_^������������VW�|$��tHh w���
P����t8�t$��t0h w����O����t ;�t������W���Z��W�������_�^�_2�^����������j�hH�d�    PQSVW�  3�P�D$d�    �ى\$3�9{�s�|$�%t�F;�tWP���%�~�~�~���D$�����I����L$d�    Y_^[���������V��F�V����;�uJ��   v��|�nf ;�}�������   ��;�}8P���G����N����F���N^�N�����F����V��R������N����F���N^����V��������D$t	V諃������^� ��j�hx�d�    PQV�  3�P�D$d�    ��t$�D$�T�H�N�P�V3ҍN�$Y��P�T$��T�Q�Q�Q�����ƋL$d�    Y^��� ������V��������D$t	V��������^� ��j�h��d�    PQV�  3�P�D$d�    ��t$�D$�T�H�N�P�V3ҍN�tY��P�T$��T�Q�Q�Q�����ƋL$d�    Y^��� �����̃�SUV3�W���l$�l$�����9o�wt�F;�t�UP�B���Љn�n�n�\$$�L$Q�T$�G Rh � @�ˉD$(�(肶����u_^]2�[��� �|$�D$$ ��   �D$P�ˉl$��k������   �D$9G}P�������D$��~%�S���x������������t��;l$|��;l$|Y�L$Q���D$    �k����tA�D$��~$P���$-���l$U����(���WU���lk����t�T$R���Lk����t�D$$��輩�����&����D$$_^][��� ������j�h��d�    PQV�  3�P�D$d�    ��j������D$���D$    tV���J����L$d�    Y^���3��L$d�    Y^���������j�h�d�    PQV�  3�P�D$d�    ��j�~�����D$���D$    tV���z����L$d�    Y^���3��L$d�    Y^���������S�\$��UVW��}S3�9n�  �~��x"��k�d���$    �N��F�������d;�}�N��PUQ����_�n�n�n^][� �F;���   �N��PSQ����3�;ŉF��   �N��+�k�dk�dR�UQ�� �F��;�};�ȋ�k�d+п%�F�t� `T�h�h�h�x�h�h�h�h ��d��u�_�^^][� ~M���;�|��+�k�d����N��s�����d��u�9^~�^�N��PSQ�Ή^��3�;ŉFu�n�n_^][� ������������j ��T�������U�l$V��;�tX�ES3�;��^[��^]� 9F}P�t���9^t�E;ÉF~�W3����E�N�P��0�������d;^|�_[��^]� ��^]� �����V��j ��T� ����D$t	V�c~������^� ���������̋��@   �@����� �Y3��@�T�H�H�H��������j�hC�d�    PQVW�  3�P�D$d�    ��t$��Y�~j ���D$   ����j ���D$ ��T�y����T�L$d�    Y_^����V��L$�FP�����F^� ��������̋L$���3����  �$� �j�p{�������  ���>���j�W{��������   ���U���j�>{��������   ���l���j�%{��������   ������j�{��������   ���j���j��z��������   ������j��z������tp������j��z������t[������j�z������tF���2���j�z������t1���=���j�z������t������j�qz������t������3������4�M�f�������������������������̃�,UVW���|$�/����t$<�D$(P�L$Q3�h � @�Ήl$�l$4�K�����u_^3�]��,� �|$S�Ä���  �W R����g���؄���  �GP���e���؄���  �OQ���g���؄���  UV�OH�%���؄���  V�O0��.���؄��{  �T$0R�D$Ph � @�Ήl$$�l$<觯���؄��S  �|$�l$@�Ä�t�L$@Q���e���؄�t�T$@R�O`�����9l$@�l$(��   ����   �D$4P�L$ Qh � @�Ήl$(�l$@�:����؄���   �|$�Ä�t{�T$ R�Ήl$$�d���؄�te�D$$P�Ήl$(�d���؄�tO�L$ Q���������;��|$8t4�T$$�W��PV���Ҋ؄�u��j������L$�D$8P��`�m}���|$��貢����u2ۋD$(��;D$@�D$(�'�����萢����u2��.��t*�|$,|#�L$@Q�Ήl$D��c���؄�t3҃|$@�W���S�����u2���[_^]��,� V��N�V;�uL��k�d=   v��|��z ;�}�������   ~�	;�}UP���:����N��k�dF���N^�k�dN�����Fk�dFt$3�� `T�H�H�H�@%�H�H�H�H �N��k�dF���N^�����������V��������D$t	V�y������^� ��j�hh�d�    PQV�  3�P�D$d�    ��t$�D$�T�H�N�P�V3ҍN��Y��P�T$��T�Q�Q�Q�����ƋL$d�    Y^��� �����̃�UVW�q3�W�������l$�D$P�L$Qh � @�͉|$�|$諬����u	_^]��� S�T$R�͉|$ �b���؄�tB�D$9F}P��������D$��~)U���6�����������t��;|$|��j ������2ۋ��N�����u2ۊ�[_^]��� ������������j�h��d�    PQV�  3�P�D$d�    ��j�u�����D$���D$    tV���z����L$d�    Y^���3��L$d�    Y^��������̸x�����������VW�|$W���"�����   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   �P���   �H���   �P_���   ��^� ������������������� ��������SV�t$Wj j��h � @������؄�t$���   P���cs���؄�t���   W��蟖���؋��F�����u	_^��[� _^��[� ��SU�l$3�V�D$�D$��D$P�L$Qh � @��脪���|$��t2���W���T$���   �$���������t�Ƹ   V����a���؄�t
W����a���؋��F�����_u^]��[��� ^]��[��� ��������̋D$h�ZP�x�����   � ������VW�|$j��j���-v������tH������$��q������t2�FP��腕������t �NQ���s�������t��(V����t����_^� ��������̸ y�����������j�h��d�    P��xSVW�  3�P��$�   d�    ��3�9F������u6��$�   ��th [P�qq�����ǋ�$�   d�    Y_^[�Ą   � �N���$�   �BS�Ћ���u��t�h[S뷍L$X�(��j �L$\Q�NǄ$�       ��� �T$R�L$\輊���x�D$(P�L$\�[)���@�����Dz!�L$@Q�L$\葊�����X����Dz�   �3���th�ZS�p�����L$XǄ$�   ������(����� ����6��������������th�ZS�lp����3�������̃�SV��NW3�;ω>t	��Pj�ҋ\$�D$P�L$Q�ˉ~�|$�|$�Dt���|$����   ;ǉ|$t�T$R���B]����;�tl�D$+�t��t_^3�[��� �   ��>�D$P�ˉ|$ �)?���؋D$;�t.P�[����;ǉFu�L$3�;�t	��Bj��_��^[��� ��_^[��� �����̸�y����������̸   ����������̋��   ���������̋D$���   � ��̃�P��V�L$ �N�T$$�V�L$(�N�T$,�V�L$0��T$4�P�L$�H�T$�P�L$�H�T$�P�L$�L$ �T$������L$������D$TVP�L$@Q��������L$8�����T$R�L$$�o����$��4������z�����P���[����z
��$��PÍD$8P�L$�0����$��P�o� ����̃�V�t$ j ���o������������z%j���W������������zVh��D$P�Vh(��L$Q�+�����L$0��P�Q�P�Q�P�Q�P�Q�@���A^����������������VW�|$��t5hx����;����t%�t$��thx����;����tW������_�^�_2�^�������������j�h��d�    P��VW�  3�P�D$ d�    ��t$������   ���D$(    �LZ������D$P�x��8�����N�P�V�H�N�P�V� 0�F�0�N�0�V �0�F$�F(   �`/���   �d/���   �h/���   �l/�����   �T$���$������ƋL$ d�    Y_^�� �V���LZ����D$t	V��o������^� �����������̃���SUV��W����n�T$���$��������\$��N�$�L$(�e����F,�^(3�;�t�K���QWP蘭 ���T$�{�|$�|$�|$ R�D$P���p���|$��u@��t<V���Y������t-U���[������t�L$Q����Z������tS����`����_^][��� �V�t$��th y���9����t��^�3�^����������������U������4SV��F ��W�t$,|����|�   ���   t";�t,��t�]��th�[S�k����3���]����   ��]�F0���D$(}��th�[S��j����3�_^[��]� 3�����   �53ۋv,��������Aza�H+�����AuR���T$�L$@�$�����P�N������t4�5�V����D{"��4�^ ����z����8;|$(})�t$,��؋E��tWh�[P�=j����3�_^[��]� �ظ   _^[��]� ���������������SVW�|$j��j����m����3�;���   �FP���$h����;���   �N Q���h����;�t{�VR���k����;�ti�F$P���k����;�tW�~ Uu=�n0;�l$}�\$��U����g��;���~3��t)�N,�W�+�������8;\$|��t��V���i����]_^[� ������V�t$��th�y���k7����t��^�3�^����������������W���O腯������u�D$��th@\P��h����3�_� SU���   V3���~&�\$���   �<� ��t�S�������t/��;�|�^][�   _� ��t+Vh,\S�h����^][3�_� ��tVh\S�uh����^][3�_� ���������QUV�t$Wj��j���Kl����3�;���   �EP���C�����;���   ݅�   �����$��g����;���   ݅�   �����$��g����;���   ���   Q���f����;ǉD$tpS���   ;߉\$}�|$��S����e������~G��tC���   ��jj���k������t�P����e������t�KQ���4������;|$|��D$[_^]Y� �����������́�   W����$�   3���|];��   }U���   ���I��tE��BdV�Ћ���t6��Btj���ЍL$��_����WhhY�L$�.}����RD�D$P���ҋ�^_�Ā   � ���QSU�鋅�   VW�D$�   3�;\$}CS���Z�������t.�۸   u�D$ �L$��R8P�D$ PQ���ҋ���Pj���҃���u���_^][Y� �����V��~ ��[t%�F��tj P��[�F    �F    �F    ^�����������V��~ ��[t%�F��tj P��[�F    �F    �F    �D$t	V�/i������^� ������j�h+�d�    PQ�  3�P�D$d�    h�   ��f�����D$���D$    t�������L$d�    Y���3��L$d�    Y������������j�h[�d�    PQVW�  3�P�D$d�    ��h�   �f�����D$���D$    t���������3����D$����tW�������ƋL$d�    Y_^��������������V������T$�N�$��������\$��N�$�����3��F,�F0�F4�F(%��^������������U������4S���V���W�}���\$��$h�\W�`d��hx\W�Ud���� �CP����f��hl\W�<d�����KQ���g���C0PhX\W�D$H�d��3���9t$<~I��|;s0}�S,�������$hT\W��c���D$L�����;�}h�fW��c������;t$<|�h�&W�c����_^[��]� V�t$Wh]V���c���G ���� t��t��uh]�h�\�h�\V�oc����h�&V�ac�����O��a����u��7Php,V�Ac�����O$��a����u��7Ph�\V�!c����� u=U�o0Uh�\V�c������~S3ۋO,V��c�����8��u�[h�&V��b����]_^� ������j�h��d�    PQVW�  3�P�D$d�    ��t$�2� 3��N�|$�4]������ݞ�   ����ݞ�   ǆ�   �[���   ���   ���   ǆ�   �����L$d�    Y_^�������j�h��d�    PQSUVW�  3�P�D$d�    ��t$�4]���   3�3�;��D$    ~?���$    ���   �<�;���t��O;�t	��Bj��W�e������;��   |�9��   ���   �D$ ��[t�G;�tSP����[�_�_�_�N�\$ ������D$ �����\ �L$d�    Y_^][�����������j�h��d�    P��SVW�  3�P�D$$d�    �ً��   W�L$舉��3�;��t$,~!V�������D$�D$P�L$�dg����;�|ߋL$<�T$8�D$4QRP�L$ �%� �L$���D$,�����b����ËL$$d�    Y_^[�� � �����������U������xS�_V�L$8�\$4�����D$8P�sHV����V�C�t$D�*����T$D��������;����Auo�KH��Q�����$����3�9��   ~@��|;��   }���   ���3��D$8�Hh�=h(����$�� ��;��   |�݇�   �D$8ݟ�   ��؍L$P�h�����=�D$XP�L$TQ��=���ĉ� >�H�>�P�>�H�>�P�H��轣���D$P������;���������D$X{(����������At�D$`����������At����^[��]��������\$�L$H���$�o���3�9��   ~E��|;��   }���   ���3��X�D$8P�L$l�k����L$hQ���O� ��;��   |��\$4�D$X���\$�T$x�D$`���$R�ҡ�����P�S�H�K�P�S�H�K�P^�S[��]�����������U����j�h+�d�    P��  SVW�  3�P��$  d�    �ًuj ���`^�����%�$���5����A��  �s�    ��$�   �uV��$�   Ǆ$$      �٧����$  ��V����$�  ��V���L$��V���CPhhY��$  �t��hhY��$�   P��$�  ��s����$  Q��$  RV��$�  P��$�  ��W������W����    �|$�j �L$�W��j ��L$�X�W����j�L$�X�W����j�X�L$�vW����j�X�L$�fW����j�X�L$�VW����j��L$�GW����j�X�L$�7W�����Xj�L$�'W����j�X�L$�W����j�X�L$�W����j��L$��V����3��X9��   ~,���$    ���   ���J��@D�T$R�Ѓ�;��   |ݍ�$�   Ǆ$   ��������uV�K�:����ȋ��L$����V���D)���D$��$  d�    Y_^[��]� �������̡�=� >��(S�مۋ�=V�t$4��>�N�>�V�>�F�N�VttW�D$P�x�~'��P���(������tUhx���*����tE݇�   ��݇�   �L$,�\$�$Q�K譞����H��P�N�H�V�P�@�N�V�F_��^[��(� V��F�V;�u=��    ��   v��|�  ;�}�������   ��;�}P���f?���V�F��    �N�V�����N^���������j�h[�d�    PQ�  3�P�D$d�    h�   �%\�����D$���D$    t��������L$d�    Y���3��L$d�    Y������������V���H����D$t	V��]������^� ��j�h��d�    PSUVW�  3�P�D$d�    ��\$$;��  ���   3���~:���   �4�����t�     �N��t	��Bj��V�V]������;��   |ƃ��    |
ǅ�       S���w �s�}�    󥋋�   ���   ���   ݃�   ݝ�   ݃�   ݝ�   ���   9A}P��=��3�9��   ~kj��Z�������t$$3�;�L$t(���   ��� ���N9Ht�@��ȋBd�ЉF�3��L$$Q���   �D$ �����t$(�_����;��   |��ŋL$d�    Y_^][��� ��������U������4SVW�}�񋆨   Phd^W��X��݆�   ���$hL^W��X��݆�   ���$h8^W�X�����L$(Q���p����D$8���\$�D$H�\$�D$@�$h ^W�{X���F���\$�F�\$�F�$h^W�YX���F0���\$�F(�\$�F �$h�]W�7X���FH���\$�F@�\$�F8�$h�]W�X���F`���\$�FX�\$�FP�$h�]W��W�����   S�\$Hh�]W��W����,���D$     ~s���   �D$ ���; uhp[W�W�����;uh\[W�W�����{ uhD[W�W�����h8[W�zW���K��B��W�ЋD$ ��;D$$�D$ |�_^[��]� �̃�SUVW��h(��^h�=��賛���荮�   �] ��   ��D$���   ���   �D$� �����G3�;�t�O��QVP�|� ���L$$�T$R�D$P�w�t$�t$ ��Z���|$����   ����   �L$$S�+E����3�;���   U�l$(���bD����;���   �L$Q���KD����;���   �T$R���C����;���   �G;�t�O��QSP�ӗ ���T$$R�͉_�\$(�mC����;�t]�D$$;�~UP���V:���\$���D$;D$$}=������j���FW����;�t��X�3�;ÉtU���x������3��D$;�u�_��^][��� �������������U����j�h��d�    P��dSUVW�  3�P�D$xd�    ��E���D$8��   �<�    +����3ۋE�9X4�p(�%t�F;�tSP���%�^�^�^�Ej8�SP赖 �u����t$<�t$@��$�   t<�����N�T$�$�6�������\$��N�$� ����F(%�^,�^0�^4�D$8����8;�Ǆ$�   �����D$8�O����]�L$xd�    Y_^][��]��E    �L$xd�    Y_^][��]��������������j�h��d�    PQVW�  3�P�D$d�    ��h�   �U�����D$���D$    t���W������3����D$����tW�������ƋL$d�    Y_^������������VW�|$��t5h�y���"����t%�t$��th�y���"����tW���F���_�^�_2�^�������������W���G�W;�uG��    +���Ɂ�   v��|�Q�$ ;�}�������   ��;�}jP���޷���`��    +ЋG�|�4 V�t�(�%t'�F��t j P���%�F    �F    �F    �G�W��    +ȍ�P���]1��^�O�G��    +у��O��_���V��j ��[�P����D$t	V�V������^� ����������VW�|$��t5h y���� ����t%�t$��th y��� ����tW������_�^�_2�^�������������j�h#�d�    PQVW�  3�P�D$d�    ��t$���3��N�|$��^�F�����7O���`/�F�d/�N�h/�V�l/�N$�D$�F�~ �O���F(�[�~,�~0�~4�ƋL$d�    Y_^����j�h^�d�    PQV�  3�P�D$d�    ��t$��^�N(j �D$   ��[������N$�D$�M���N�D$ �M�����D$������$���L$d�    Y^��Ã�SUVW��3��G�����o�E �E�E3��E�O�w �M���O$�M���O(�L$�>����\$$�D$P�L$Q�ˉt$�t$$��T���|$���  ��t�GP����=�������D$    ��   �T$R����=��������   �D$�� t#��t��t3��   �G    ��G    ��G     �GP���|B������tu�G$P���jB������tc� u]�|$���r����D$$P���D$(    �N=������t7�D$$��~/P��致��3���I ;|$$}�L$�A���S���y���������u��|$|U���!?��_^]��[��� _��^][��� ��������j�h��d�    PQ�  3�P�D$d�    j8��P�����D$���D$    t�������L$d�    Y���3��L$d�    Y���������������j�h��d�    PQVW�  3�P�D$d�    ��j8�TP�����D$���D$    t���������3����D$����tW�������ƋL$d�    Y_^���������������V��������D$t	V��Q������^� �̸�z�����������j�h��d�    PQV�  3�P�D$d�    ��t$�3���N�D$    �`_�mK��3��F�����F�F�F�F�ƋL$d�    Y^��������j�h�d�    PQV�  3�P�D$d�    ��t$�`_�N�D$    �"J�����D$�����s!���L$d�    Y^�����VW�|$j��j���Q������t2�FP����K������t �NQ���iO������t��V���M����_^� ��������������̃�SUV��W�^�~���������I���l$3�����F�F�F�D$�D$�D$P�L$Q���'Q���|$��u>��tW���1:������tS���?�����|$|��tV���,<��_^]��[��� 3�_^][��� ���j�hK�d�    PQ�  3�P�D$d�    j ��M�����D$���D$    t��������L$d�    Y���3��L$d�    Y���������������V�t$��th�z���k����t��^�3�^����������������j�h{�d�    PQVW�  3�P�D$d�    ��j �4M�����D$���D$    t���J������3����D$����t4W����$���GP�N�O���O�G�N��V�H�N�P�V�@�F�ƋL$d�    Y_^���VW�|$��t5h�z�������t%�t$��th�z�������tW���&��_�^�_2�^�������������V�������D$t	V�[N������^� ��VW���O�I������u��7�G�|$Ph�_W��J��Vh�_W��J����_^� ��V�t$��th�{��������t��^�3�^���������������̸�{�����������V��W�|$���O�N�W�V�G�F�O�N�W�V�G�F�O �N �W$�V$�G(�F(�O)�N)�W*�V*�G+�F+�V,�R�N,�G,P�ҋF<�@�N<�W<R���OL_�NL��^� ��������������D$W��������������A��   ���L$����|$������������+������������������   ������_�h������������������D$�����_~v������+���������������������������_~Z������tP������3��_� �D$�م���|4�|$�L �����?3��_� ��_����������� ��������������_� ��������U�������   S�]��	VW��~�C��P�+d�������|$<�
�L$`�L$<���E�T��f�T$D��������Az�   �3��D�(�����E�f ��������u�   �3��~�D�8�T$X�������T$Pu!W��S�ك��\$���$�C����D$X�D$P�,�����~ ���_~�K�����t������3������Ƀ~uR��S���\$���$������(���~ ���Z~����zt�ˁ�����3�����3�9]�\$P��   �D$<����D$@�E�K3����\$H�L$L|f�|$L�L$@���|$X����+߉\$H�\$X�A�� �NH�� �� ���J��X��A(�NH�J��X��A �NH�J��X��A�NH�J��X�uT$D�\$P;�(�T$H�L$<�ыT$D����NH����;��L���X�~�\$L�D$@;]�\$P�F���_^[��]� ��������VW�|$��;~tkS3�;�~J9~~�~�N��PWQ����;ÉFt@�V;�~��+ʍ�����Q���SR�� ��[�~_^� �F;�t�SP�B�Љ^�^�^[_^� ���SW�|$����~eU�l$��|[V�t$��|Q;�tM�C�/;�C;�?�K�>;�~�;�}��P���6����C����R�L� �������Q�R�� ��^]_[� ����������V��~ ��_t%�F��tj P�`�F    �F    �F    ^�����������VW�|$��;�tD�G��_�F    ��^� 9F}P�Tm���N��t�G�F�W�����PRQ�� ��_��^� ���������V��~ �`t%�F��tj P�`�F    �F    �F    ^�����������VW�|$��;�tA�G��_�F    ��^� 9F}P������N��t�G�F�W����PRQ�F� ��_��^� ������������V��L$��|6�F;�}/+���P�APQ�������F��F����NjPj Q�� ��^� ����������̋D$�L$����PQ��_����� �����V��~ ��_t%�F��tj P�`�F    �F    �F    �D$t	V�/G������^� ������V��~ �`t%�F��tj P�`�F    �F    �F    �D$t	V��F������^� �����̋D$SU�l$j UP���;�  �Ѕ҉T$��   ��V�sLW3���|t�KH�V�����8���<�    �A���������Au��������������Au������A(��������Au������AP��������Au����؁��   ��u��T$;�}'�CH���L�+����������Au����؃�(��u�D$����_^t� ����@���X�@���X���t�E ���] �E���]�E�]][� ��][� ������j�h��d�    PQSVW�  3�P�D$d�    ��t$h@h`�jj�~W��� 3ۉ\$�F,�_�^0�^4�^8�F<`�^@�^D�^H���D$��^(�^)�^*�^+�����N����9^H��|�^D�^L�L$d�    Y_^[����������j�h�d�    PQSUVW�  3�P�D$d�    ��t$3ۍn���D$    ��^(�^)�^*�^+�#����N����9^H�~<|�_�^L9_�D$ �`t�G;�tSP���`�_�_�_��,9^�\$ ��_t�F;�tSP���`�^�^�^h@jjU�D$0�����R� �L$d�    Y_^][���������������j�hH�d�    PQV�  3�P�D$d�    ��t$�s  3��N�D$�$`�F�����ƋL$d�    Y^�����������̃�SUV��3�W�~�ω�^(�^)�^*�^+������n������9^H|�^D�L$$;ˈ^L���   ��@lS�T$R�Ћ��P�W�H�O�P�L$�W�������@lj�T$R�Ћ�M �P�U�H�M�P�L$�U��������7�����t���,�����t_^]�[��� �ω�^(�^)�^*�^+�G������@���9^H|�^D_�^L^]��[��� _^]2�[��� �������������V��F�V;�u<������   v��|��� ;�}�������   ��;�}P���7����F����VjPj R聀 �N����F�����N^�����������j�h{�d�    PQ�  3�P�D$d�    jh��?�����D$���D$    t��������L$d�    Y���3��L$d�    Y���������������j�h��d�    PQVW�  3�P�D$d�    ��t$�$`�~j ���D$   �����N��t;�t	��Pj�ҋ��F    �D$ �F������D$�����  �L$d�    Y_^��������VW�|$��;�t\�N��t;�t	��Pj���F    � t���  P�ΉF�a  �W���  S�^��W�������������P���	���[_��^� �U����j�h��d�    P��$  SUVW�  3�P��$8  d�    �ًs43��{L �t$(��  9;��  ;���  ��$�   �L7��9{H�K<��$@  |�y9q}V����;���  �D$(�D$     �D$$��$    �K<�h����s0t$ �
   �|$\�sj �΋������j�D$`��� �\$8����� �d$\�T$<�D$4������������Dz�������\$4���������Dz���\$<��؍{j ��蛥���D$d� j���\$H舥��� �D$d�����T$�D$D������������Dz�������T$D���������Dz�������T$�����D$\�   �U �E�]�E���U�] �0'�D$4���](���D$<���]0�������]8�������]@���]H�\$t������  ��$�   �	�����$�   �������$�   �����D$dj j ��$�   Q���$�   R��$�   P���\$݄$�   �$�YP  ����  �D$<�D$4������Au������\$,�D$�D$D������Au����؍�$�   �\$L菲����;������z�|$t�D$,������Au�\$,��؍�$�   �[�����;������z�|$t�D$L������Au���
���D$L��ـ{( t�D$D������Au�����{) t�D$<�D$,������z����D$,���ɀ{* t�D$������Au����܀{+ t�D$4������Au������0'�������](���������]0�����]8��  �sj ���?���� �\$\����D��   �Ej ���\$����� �\$����D��   �{) u;�{+ u5j���E   ����� ���]赣���=0'���](襣���=0'�]0�{( �@  �{* �6  j���E   訢��� ���] �l����=0'���]8�\����=0'��  �E j���\$�q���� �\$����Dzd�Ej ���\$�T���� �\$����DzG�{) �q����{+ �g���j ���E   �#���� ���]����������](�٢�������1����E j���\$����� �\$����D��   �Ej���\$�ϡ��� �\$����D��   �{) u7�{+ u1j ���E   袡��� ���]�f���������](�X��������]0�{( ��   �{* ��   j ���E   �]���� ���] �!���������]8�����   �E j ���\$�.���� �\$����D��   �Ej���\$����� �\$����Dz~�{) u;�{+ u5j������� ���]诡���=0'���](蟡���=0'�E   �]0�{( u7�{* u1j ��誠��� ���] �n���������]8�`����E   �����]@�D$ (�l$$�R����t$(VV��$�   � � ����QƄ$D  �]R������3���D$$�T$,��   3��D$4�D$ �C@D$ �L$4� �T$$�\$L3��@�C0�\$T3��D���D$T�K@�D$Pj ���\$��D$d�$����U��$�   衑 �D$������P;t$(|��D$ P�D$4(��;l$(|��t$$��;j V����$�   �$�<� �|$(;��l$,u#��;UVW����$�   �$�� ��t�CL�{L ��   3���|Y�W���3Ƀ��E�4�    ��$    �k@�@��\)H�k@�@��� ݜ)�   �k@�@���@  ���\)��@�k@�\)�uǋl$,;�}$�������$    �D� �K@�\H����P;�|�T$$R�Q������$�   Ƅ$@   芕 ��$�   Ǆ$@  �����S1���CL��$8  d�    Y_^][��]����������j�h�d�    PQVW�  3�P�D$d�    ��jh�46�����D$���D$    t���
������3����D$����tW��������ƋL$d�    Y_^���������������VW�|$��t5h�{�������t%�t$��th�{�������tW������_�^�_2�^�������������V��������D$t	V�{7������^� ��U�������   SV��M�A�����+�����W�t$P~�}�ˁ�����3����|������D$G�  ��~��    P�.O�����D$K���t$L�
�L$X�L$L��T$P�JD����   �D$H    �L$T�E�E�L$P�I@L$HVP���\$�E�$����3���|R�E�S��N+u�������<�    ���A�� �@؃� ���X��D��@��X��A��@��X��@��A��X�uЋt$L;�}�M�֍�+ы�+�������@��X�u�D$HP�l$T�O����D$G�T$X;�tV�wN���D$K��_^[��]� �������U������  S�]V�u W�L$4��$�   �D$0   ���������l$0y�E��}��$�   �   ����˃��   �U(�ER�U$RWQ�L$DP���\$�E�$�  ;��ЉT$0tn݄$�   �M���݄$�   �^݄$�   �^��   ݄$�   ������݄$�   ��\�݄$�   �\�݄$�   �݄$�   �X݄$�   �X�rV��$�   ������Q��$�   �ڦ�������R��$�   �Ʀ���[��Q��$�   賦�������R��$�   蟦������Q��$  茦���M�T$0����  ��~!�A�����+������P�L���������$  �U�E�L$4WR���\$���E�$����������D$0�F  �L$@�g����D$@P��$  Q��$�   R��$�   P�E$��$�   Q��$�   RP�q� �D$\����} ���D$H��F�^�D$P��F�^��   �L$p������L$X�����L$XQ�T$tR��$  P��$�   Q��$�   R��$�   P��$�   Q�ٯ �G�D$\�����D$p����������G�D$H���D$x������D��\��G�D$P��݄$�   ������D��\����G����D$X��������O�D$`����F�^�O�D$h����F�^��$  ;�t	W�9K�����D$0_^[��]�$ _^��[��]�$ ��������������V�t$��th�|��������t��^�3�^���������������̸�|�����������V���7  3��F�F�<a��^�������V���7  �D$�F�<a�F ��^� ��K������������V��~ t"�N��T$�@R�Ѓ�VjP蜈 ��^� �D$��VjP腈 ��^� ��������������VW�|$��;�tW�~L  �G�F�O�N_��^� ������������<a�A    �7  ��������������V���F    �A���D$;�u3��F�F^� �F �F^� ��V��N3���t!W�~����~ ��t��t����   ���ҋ�_^�̃y t
�I��@��3�� �����������VW�|$��FPhbW�-�����~ t�N��BW��_^� �y t
�I��P4��3���������������j�hY�d�    P��VW�  3�P�D$ d�    ���D$    �t$0���D$(    �n���� �D$(    �D$   t3�9D$4����D$4� t/�O��RlP�D$P�ҋ��P�V�H�N�P�L$�V������ƋL$ d�    Y_^�� � ��������������3�9At78At�D$�I�T$V�1P�FpR��^� �D$�I�T$V�1P�FpR��^� �L$���t��L$��t�� ��� ���̀y t3�9D$����D$�y t�I��D$�Bt��3�� �̀y t3�9D$����D$�y t�I�V�t$VP�Bx��^� 3�� ����������̀y t3�9D$����D$�y t�I��D$���   ��3�� ��������������̀y t3�9D$����D$�y t'�I�D$�V�t$V�t$V���$P���   ��^� 3�� ��������̀y t3�9D$����D$�y t�I��D$���   ��3�� ��������������̋D$VW��3�� t��ȋBd�Ћ���BPjj ���ЋƋO�|$�WP���   �Ѕ�����   �G���w~�$��$��Bj�ο   �Ћ�_^� ��B�   W���Ћ�_^� ��Bj�ο   �Ћ�_^� ��Bj�ο   �Ћ�_^� ��Bj�ο   �Ћ�_^� �   ��Bj���Ћ�_^� �f$}$�$�$�$�$��������j�h��d�    P��   SVW�  3�P��$�   d�    ����$�   �^j ���ߟ�����$j���П�����L$ �$����P�L$4����j ��讟�����$j��蟟�����L$0�$谧��P�L$L�֞���D$0P�L$LQ�L$h�#���� Ǆ$�       t�t$`�O����   V�Ѐ ��t7�F���w/�$�P&�   �!�   ��   ��   ��   ��   �L$`Ǆ$�   ���������Ƌ�$�   d�    Y_^[�Č   � �%�%&&&&��������W��3�9Gt9�O�D$����   S�\$V���$S�ҋ���t� t��t	���p����^[_� ��������̀y t3�9D$����D$�y t�I��D$���   ��3�� ���������������2��y ta�T$��wX8At	�   +�����D$0�IV�t$(����\$�D$<�$V�t$8�D$,V�t$8V�t$(���\$�D$<�$VP���   ��^�4 ���̀y �D$t#��w�$��'�   ��   �	�   �3��y t�I��D$���   ��3�� �I �'�'�'�'����V���X���~ ���F�   ^�������̃y �te�y t
�D$�D$��D$�D$�D$<�T$�I����   ��(�\$ �D$\�\$�D$T�\$�D$L�\$�D$D�$R�T$0�Ƀ��\$�$R���@ �y t
�D$�D$��D$�D$�y t5�T$$�ɋI����   R�T$$R�T$$R�T$$R�T$$R���\$�$���$ ��3����$ ����3�8At�   +T$��T$9At��w�I�D$����$R���   ��� �����V��~ t8�N�D$����   W�|$���$W�҅�t�~ t����   ����_^� 3�^� ��������̃y u3�ËI����   ������������2��y tW8A�It)�T$�D$����   R�T$R���\$�D$$�$��� �D$�D$����   P�D$P���\$�D$�$��� ��������������2��y tW8A�It)�T$�D$����   R�T$R���\$�D$$�$��� �D$�D$����   P�D$P���\$�D$�$��� ��������������j�h��d�    PQV�  3�P�D$d�    j��%�������t$���D$    t+���-  �<a�F    �F �ƋL$d�    Y^���3��L$d�    Y^�������j�h��d�    PQVW�  3�P�D$d�    ��j�d%�������t$���D$    t���,  �<a�F    �F �3����D$����t;�tW����A  �G�F�O�N�ƋL$d�    Y_^��������������VW�|$��tEh�|���������t5�t$��t-h�|��������t;�tW���rA  �G�F�O�N_�^�_2�^�������������V���<a�F    ��+  �D$t	V�n&������^� ����̸�}�����������V�t$��th�~���+�����t��^�3�^���������������̸�~�����������SU�l$V��W�    �������   �P���   ��������   ���   ���   ���   ���   ���   ���   _���   ���   ^]���   ��[� ����j�h;�d�    PQV�  3�P�D$d�    ��t$�*  �N�D$    �\b�d��h@h`�jj���   P�D$(�Ê h@h`�jj���   Q�D$(褊 �ƋL$d�    Y^���������������SU�l$��;���   VWU�?  �u�{�    󥋅�   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ����   �P���   �H���   �P_���   ^]��[� ����������+���   ������V��L$�FPh�   Q�z ���   Rj P�{z �ƨ   Vj P�lz ��$^� �������SV�t$��W���\$�{��    ��$���   ��肛�����荻�   �\$�����$�g�����N�V���   �F���   ����   �O���   �W���   �G���   _���   ^���   ��[� ���������j�h��d�    PQV�  3�P�D$d�    ��t$�\bh@jj���   P�D$$   ��� h@jj���   Q�D$$�݇ �N�D$ �������D$�����(  �L$d�    Y^�����������������V��N�e����tE���   薉����t6���   臉����t'���   �x�����t���   �i�����t	���^� 2���^� ��̋D$h0cP������� �����������VW�|$j��j���"������tb�FP���@������tP���   Q����A������t;���   R����A������t&���   P����A������t�Ƹ   V���A����_^� ��������������̃�S�\$V��D$P�L$Q���D$    �D$    �"��������   �|$��   �VR���S������t&���   P���������t���   Q���������|$���   ���   ���   ���   �Q���   �Q���   �Q���   ���   ���   W���   �W���   �W���   �W|��tQ���������tW���y����_^[��� �������������U������   SVW�}W����������   j �^8�L$4�B����D$ �F ���   j �D$<�L$8�&����L$ �S����$�   �$R�D$8���Տ���L$H�T$8���P�D$\PQ����$�   �$P讏����P��$�   Q���ˎ�����Ď���L$0j蹅���L$4j�D$,誅���T$(�S�D$$����$�   �$P�\����T$H��P�D$$� �L$DQR����$�   �$Q�5�����P��$�   R���R������K���W���e�����Ä���  j ���������%�$����4����A�n  �D$XP�L$|Q��������T$X�H�L$\�P�T$`�H�L$d�P�T$h�@�L$@Q�T$|R�ωD$t�����L$@�P�T$D�H�L$H�P�T$L�H�L$P�P�D$ P�L$tQ�L$d�T$\�T$`���ĉ��$�   �H��$�   �P��$�   �H��$�   �P�H��2��!_������   �L$@�T$(R�T$H�D$<P���ĉ�L$h�P�T$l�H�L$p�P�T$t�H�ΉP��^����tb�D$8�D$p������zM�D$(�\$ ����Au>�L$4�Ƀ��\$�$豕���D$(�L$0���\$�D$0�$薕�����_^[��]� ����_^��[��]� ��������Q�|$ �$    t���   ����   �D$���Q�P�Q�I�P�HY� �����j�h��d�    P��V�  3�P�D$d�    �T$(��@lR�T$R�ЍL$�D$     �
����t$,�L$��k����^�L$�����L$���D$ ���������ƋL$d�    Y^��� �������D$3�9D$V�������   �D$�L$PQ���$j��蟂�����$j ��萂�����$�5� �� ^� ��������������W�|$���   tV�q�    �^_� ���D$0�D$$�T$ ���\$�D$8�$P�D$0�D$(R�T$ P�D$ ���\$�D$8�$RP��6  �4 �����������S�\$��V��wI����W�<0���   菅�����   脅����_�N8u�N �$����NP�����N��[��^�   [� ^3�[� ��̰�@ ����������̃�SV��W�N�_�����   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   �L$���   �L$�D$�T$�|$���   ���   �g���_^�   [��������������U������4��SV�T$���\$W���   ���   W��脖����t:�E�����$蠀�������$�S����]��������\$�������|$�\$���   ���   W���2�����t:�E�����$�N��������$�����]��觀���\$ ��蜀���|$ �\$ �E���\$�D$8�E�N�$P�WY���D$(�M �]��D$0�U�Y�<�    �D$8�Yσ�|f�F �D$������F(���Y�N0�Yσ��F8�D$ ������F@���Y�NH�Y~)�B���+������Í�   R�j W�IW ��_^�   [��]�$ ��������U����j�h�d�    P��   SVW�  3�P��$�   d�    ��}3ۅ�t	����  ��Pj �҅���  �L$T�p	 ��PlW�L$0Q3ۋΉ�$�   ��S�L$0Ƅ$�   �v~��������uW� �D$L�\$�E�$P�F9  ��L$T�P�T$X�H�L$\�P�T$`�H�L$d�PW�L$0�T$l�#~��� ���\$�E�V�E�\$� �D$L�$P��8  ��L$T�P�T$X�H�L$\�P�T$`�H�L$d�Pj�L$0�T$l��}���E���\$� �D$L�$P���8  ��L$l�P�T$p�H�L$t�P�T$x�H�L$|�PjP��$�   �m�����D$(;�Ƅ$�   t�L$TQ���~�  ���3��FH   �T$,�V8�D$0�F<�L$4�N@�T$8�L$,�VD��$�   ������L$TǄ$�   ����������Ƌ�$�   d�    Y_^[��]� �Ë�$�   d�    Y_^[��]� �������������U����j�hP�d�    P��   SVW�  3�P��$�   d�    ���]���-  ��PlS�L$hQ����j �L$hǄ$�       �k|���5�����Dz8j�L$h�Q|���5�����Dz�E��P�L$d�H�T$h�P�L$l�T$p�L$T�|�������48���   ���   ���   �t$<�ƨ   �L$D�N�T$H�D$L�L$P��RlS�D$xP��Ƅ$�   ��P�EP�L$\Ƅ$�   �g����L$tƄ$�   �v����L$T�|����uPƄ$�   �L$D�X����L$TƄ$�    �G����L$dǄ$�   �����3���3���$�   d�    Y_^[��]� �|$<�ǈ   V���Ǒ����t"�L$T�T$X�D$\�L$D�L$`�T$H�D$L�L$P�ij �L$X�{��� �����$�W{�������$�
{���\$<j�L$X��z��� �����$�,{�������$��z�����\$�L$T�D$L�$舌���L$D�{����Ƅ$�   ������T$D�D$H�L$L��T$P�F�D$T�N�L$X��D$`�V�T$\�O�W�L$D�G� ����L$TƄ$�    �����L$dǄ$�   ����������   ��$�   d�    Y_^[��]� ��������������U����j�h��d�    P��   SVW�  3�P��$�   d�    ���u����  ��PlV�L$hQ���D$W �����>���   ���   ���   ���   �D$T�FǄ$�       �L$X�T$\�D$`�E��RlP�L$xQ��Ƅ$�   ��j ��Ƅ$�   �Ey���Mj �D$T�Gy���D$P��D$N����{�D$N �L$tƄ$�   ������|$N taj �L$h�D$S��x���Mj �D$T��x���L$P�j �L$X��x���Mj �D$T��x�������   �$�y�������$��x���T$P��M��@lQ�T$xR����j��Ƅ$�   �x���Mj�D$T�x���L$P��D$N����At�D$N �L$tƄ$�   �����|$N ��   j�L$h�8x���Mj�D$T�:x���T$Pj��L$X�x���Mj�D$T�x�������   �$�Zx�������$�x���D$P��������L$d�T$h�D$l���   �L$p���   �T$T���   �D$X��T$`���   �L$\�F�N�L$T�VƄ$�    �\����L$dǄ$�   �����H������$�   d�    Y_^[��]� �|$O �l����L$TƄ$�    �����L$dǄ$�   ���������2���$�   d�    Y_^[��]� ����U������4SVW����Pj �҅��D$$��   �5�W����D�T  �W �_ ����D�C  �_8�w8����D�4  ���   ��w�����!  ���   �w�����  ���   �Vw����$����A��  ���   �:w����$����A��  V�D$,SP�������L$(葄���5����A��  h�chdch�  hDc�wj�����D$$   �u�   �   j�ΉF�F    �^�^�^�^�F4�F0   ��l��Sj ���Ll��Sj���Bl�����   j ����u���N(�j���u���V(���   �Zj �u���F,j����   �u���N,�Yj ���   �}u�����$j ���nu�����T$8�$R���<0  Pj j ���Ѕ��j���   �Cu�����$j ���4u�����D$8�$P���0  Pjj ��薅��j ���   �	u�����$j����t�����L$8�$Q����/  Pj j���\���j���   ��t�����$j����t�����T$8�$R���/  Pjj���"����D$$_^[��]� �؋D$$_^[��]� �����̋�Pj ��������j�h��d�    PVW�  3�P�D$d�    ���t$���D$    ��   �L$ �>u����tt�L$ �T$$���|$0 �>�t$(�|$,���   ���   ���   ���   t���   ���   ���   ���   �L$ �D$����������L$d�    Y_^��� �L$ �D$�����e���2��L$d�    Y_^��� ���������������Q�|$ �$    t���   ����   �D$���Q�P�Q�I�P�HY� �����V��L$2҃�wB�D$�D$������z-S�Ƀ��\$����1�   �$��ӄ����������[^� ������^� ���������V�t$Wj j��h � @��������u_^� SW���F+���؄�t�G P���e	���؄�t�O0Q���1���؋��J2����u2ۊ�[_^� �����������̃�VWj83���WV�~J ���D$P�L$�|$�|$�|$Qh � @���y@����u_^��� �|$S�Ä�t,V�������؄�t�V R��������؄�t��0V���&���؋��=4����u2ۊ�[_^��� ������������SV��W�    �hY��󥍋�   袳���`/���   �d/���   �h/���   �l/_^���   ƃ�   [����������j�h�d�    PQV�  3�P�D$d�    ��t$�SJ�����   �D$    � ������D$�T����ƋL$d�    Y^����j�hH�d�    PQV�  3�P�D$d�    ��t$���   �D$    腽�����D$����膿���L$d�    Y^�������̃��  3ĉD$SV�t$(W��������D$P�L$Qh � @���D$    �D$    �>����u_^[�L$3���C ��� �|$�Ä���   �T$R���*����؄�t�|$ u-�L$�T$j���ĉ�L$0�P�T$4�H���   �P��������   P��������؄�t7W��������؄�t)���   Q��� ���؄�t�|$ ~V���   �'����؋���1����u2ۋL$$_^��[3��C ��� �̃��  3ĉD$V�t$Wjj��h � @��躥����u_^�L$3���B ��� �`/�d/�h/SU�D$�l/�L$���   �͉T$�D$�~�����~"���c�����L$�P�T$�H�L$�P�T$�D$P������؄�tA���   Q������؄�t-W���j'���؄�t���   R����-���؄�t
V���ǻ���؋��^.����u2ۋL$ ]��[_^3��B ��� �S��V���   W����������\$��{�    �$󥍋�   �������荋�   �\$���$��������\$�0'���   �$��������\$�0'���   �$����_^[����̸    �����������j�h��d�    PQV�  3�P�D$d�    ��t$��������   �D$    ��c�*������D$�����ƋL$d�    Y^��������������j�h��d�    PQV�  3�P�D$d�    ��t$��c���   �D$    �������D$����������L$d�    Y^�����������������������p  ������V��L$�FPh�   Q�Z] ���   Rj P�K] ���   Qj P�<] ���   Vh�   P�*] ��0^� ���V�t$Wj j��h � @���آ����u_3�^� Sj h � @���^����؄�t.V���@����������,����u2����tV���   �����؋���+����u2���[_^� ���̃�UVW�������t$ �D$P�L$Q3�h � @�Ήl$�l$�/:����u_^3�]��� �|$S�Ä�tc�T$R�D$(P�Ήl$,�l$ �l$$��7�����Ä�t=�|$$ � @�Ä�tV���������Ë���-����u2����tV���   ������؋��-����u2���[_^]��� ������j�h��d�    PQ�  3�P�D$d�    h�   ������D$���D$    t���K����L$d�    Y���3��L$d�    Y������������V�t$��th�}��������t��^�3�^����������������j�h�d�    PQVW�  3�P�D$d�    ��h�   �a�����D$���D$    t���������3����D$����tW���-����ƋL$d�    Y_^������������VW�|$��t5h�}���������t%�t$��th�}���������tW�������_�^�_2�^�������������j�hK�d�    PQ�  3�P�D$d�    hx  ������D$���D$    t�������L$d�    Y���3��L$d�    Y������������VW�|$��tGh�~���*�����t7�t$��t/h�~��������tW���������   W���   �����_�^�_2�^�����������V��������D$t	V��������^� ��j�h��d�    PQV�  3�P�D$d�    ��t$��  �N�D$    �\b�A��h@h`�jj���   P�D$(��g h@h`�jj���   Q�D$(��g �T$R���D$�~����ƋL$d�    Y^��� ���������U������   SVW���|$@�t$`�   �����9o������y񍏈   �D$`�L$8�D$<   ����$    �|$@�D$D���ǘ   ��0�   �D$D��T$8�L$@���\$�D$X��$P�"  ���P�V�H�N�P�V�H�N�P�V������u��D$8�l$<u��M�U3�9E��PQR�D$lPjjSj������� _^��[��]� ����������j�h��d�    P�� VW�  3�P�D$,d�    ��|$<��t.j �D$P�������D$4    �g����L$�D$4����裵���|$@��t0j�L$ Q���M������D$4   �~g����L$�D$4�����k����   �L$,d�    Y_^��,� ��U����j�hI�d�    P��   SVW�  3�P��$�   d�    ��}3ۃ��\$8��  ��PlW�L$@Q�����Ej�����$��$�   �rh�����L$<�D$7Ǆ$�   �����Ǵ��8\$7�w  W�D$hP���p����D$<��RlW�D$XP��Ǆ$�      �ҋL$<Q��Ƅ$�   �>|���L$T�D$7Ƅ$�   �i����L$dǄ$�   �����U���8\$7t�E�\$<��   ��RlW�D$XP���҉D$<W�D$hP��Ǆ$�      ������D$P�E�L$<���$Ƅ$�   �e���L$P���$�;e���L$d�\$<Ƅ$�   �ֳ���L$TǄ$�   �����³��W�L$xQ���u����D$<j�����$Ǆ$�      �'g�����L$t�D$7Ǆ$�   �����|����|$7 �+  �U���t�M;�  P�����؃����  �U���tP���������D$8��   ��u8h�   �>������D$P��Ǆ$�      t	�������3�Ǆ$�   �����؃|$8 u:h�   ��������D$P��Ǆ$�      t	���B����3�Ǆ$�   �����D$8V�������V�t$<�������E�U�G	�������ݜ1�   �1�D$<�����ݘ�   �E��0�   ��$�   d�    Y_^[��]� 3���$�   d�    Y_^[��]� ������������V��������D$t	V�+�������^� ��j�h{�d�    PQVW�  3�P�D$d�    ��hx  ��������D$���D$    t���������3����D$����tW���������   W���   �����ƋL$d�    Y_^����������j�h��d�    P��SUVW�  3�P�D$$d�    ��t$4h�dV���������~�����p  Ph�dV�����h�dV����������V���3��D$�[�|$�|$�|$ �L$Q��H  �|$0�̵��9|$~13ۍd$ �T$�P�������h�&V����������;|$|�3����.���9|$ �D$,�����D$�[t �D$;�tWP�L$��[�|$�|$ �|$h�dV�-�������`  U���|���h�&V����h�dV���������|���h0cV��������������������L$$d�    Y_^][��� ����������V�t$��th����������t��^�3�^���������������̸������������3���������������V���� �de��^��������������̋D$VP���� �de��^� ��������de� ����̸   �����������j�h��d�    P��V�  3�P�D$d�    �T$(��@lR�T$R�Ћt$,���D$     tj �L$� `��� ��t$0��tj�L$�	`��� ��L$�a���L$���D$ ����踮���ƋL$d�    Y^��� ��̋D$���t��D$��t�3�� ��3�� ��������������j�h�d�    PSUVW�  3�P�D$d�    ��l$$���D$    wE�L$(�`����t8�>j�L$,�O_��j �L$,���B_������\$��� �Gh�$U�Ѕ�t��2ۍL$(�D$���������ËL$d�    Y_^][��� ���������SU�l$V���PtWU3��ҋ�����   ��   P��������؋BxSU���Ћ���ta�L$ �D$j Q���$SWj�E� ����|>;�:�L$$��t��L$(��t*�D����\$���$�Bp��S�����_��^][� 3�S�����_��^][� _^]��[� ���j�h8�d�    P��V�  3�P�D$d�    �T$(��@lR�T$R3��ЍL$�t$ �_����t<�L$8�D$,�T$4QR���L$�$�;s�����L$ �$�r�����$�qv �� ���L$�D$ �����k����ƋL$d�    Y^��� ������U����j�h~�d�    P���   SVW�  3�P��$�   d�    �ً}���u�D$H    �v  ��Ph�L$TQ���ҋ�Ǆ$       �r�����L$\�$�g]���\$L���lr�����L$\�$�M]������4���D$L����������   ������4����   ��������A��   ������W�L$X�s���L$T�]������   �L$h���������   �L$TQ���T$t�$R��Ƅ$  �Ѕ�tm����   j �D$lP���ҍL$h��Ƅ$    �4����L$TǄ$   ���������Ƌ�$�   d�    Y_^[��]� ��������z#������Au�E����L$hƄ$    �����������؍L$TǄ$   ����萪����$�   ������P4��Ǆ$      �҃�t	����   3�W��$�   P��� ����   ����   ��$�   P���҉D$H�������   �$��]݄$�   ܤ$�   ��;������AuL݄$�   ܤ$�   �+݄$�   ܤ$�   ��;������Au݄$�   ܤ$�   �8f����u����؋���   �����$�҅�u�|$H��$�   Ǆ$   ����聩���D$H��$�   d�    Y_^[��]� �#]P]#]P]#]P]������������U����j�h��d�    P��   SVW�  3�P��$�   d�    ���u�F(3��^����D��  �F��&�PlS�L$h�\$(Q�F ���f�\$4�ҍL$d��$�   ��n���\$<�L$d�Wo���\$D��Plj�L$xQ���ҋ�L$d�P�T$h�H�L$l�P�L$t�T$p�����L$d�n���\$T�L$d�	o���T$\�D$D���D$<�����@f�����\$4���D$T���������\$L����������  ����������  �D$4�\$$����t�D$L�\$,�����d  ���L$$���L$,���������*  �����D$4�����^����uG��؋��   �؍L$Q�T$R���$j ������\$����uh�D$�^����uZ�   ��  �������AzM��ً��   �D$P�L$Q���$j ������\$����u�D$�^����u
�   �  �D$<�D$D�F��������At�����A��  ����F�����   �L$Q��$�T$R���$j ������\$�����G  �D$�^�����5  �   �+  �����D$L�����^ ����uH��ڋ��   �ٍD$P�L$Q���$j�����F�\$����Aug�D$�^ ����uY�   ��   ���^����AzK��؋��   �L$Q�T$R���$j�����F�\$����Au�D$�^ ����u�   �~�D$\�D$T�^����{�����Auc����F��F ���   �D$P��$�L$Q���$j�����F�\$����Au'�D$�^ ����u�   �����������������؍L$dǄ$�   �����s����Ë�$�   d�    Y_^[��]� ���������3�� �����������U������8VW�t$�   ���]������y��E��(�\$8��������T$X�T$`�E�\$h�L$h�T$l�T$p�T$x�E(�\$8�\$0��L$p�P�T$t�H�L$x�P�T$|�H�L$P�P�T$T�ĉ�L$X�P�T$\�H�L$`�P�T$d�H�Pt�]�����F�����@����   �E��(�\$8���E �����\$h�E(�L$h�T$l�\$8���\$0��L$p�P�T$t�H�L$x�P�T$|�H�L$P�P�T$T�ĉ�L$X�P�T$\�H�L$`�P�T$d�H�Pt�˩����@_^��]�譨����@_^��]�����U������4  SV���P4W�҃���}��W�_�0��P4����=�   �|$@���P4�������P���������E �M��S4PQW�����EP���   j ���\$���E�$�Ћ�؋B4���Ѓ�~,��E���G���X�G�X�B4��=�   ~	W�����_^��[��]� ��������������U������4  ��P4SVW�L$<����]��S���� �S�E��P�P�E ��P�X�|$@��v���P���������E(�E�L$<����   P�E$PWVj���\$�E�$����U�D$<�����������8�8�E �~9���G�[�D��Z�A�X~!�� �G�[�D��Z�A�X~	W������D$<_^[��]�$ �������������U������4  ��P4SVW�L$4����]��S�����S�E��P�P�E ��P�P�E$��P�P�E(��P�P�E,��P�X�|$@��v��P���������E4�E�L$4����   P�E0PWVj���\$�E�$����U ��D$8���E������9���v�ǍǋE$������8ǃ��D$<�E(����ǍǉD$4�E,���   ���G�E�[�D��X�E �A�X�E$�B�X�D$<�@�E(�X�D$4�@�E,�X~G���G�[�]�D��[�A�M �Y�L$<�B�U$�Z�U(�A�L$4�Z�A�X~	W�������D$8_^[��]�0 ����������U����j�h��d�    P���  SVW�  3�P��$�  d�    �ًE,�E�M(�U P�EQ�MRPQ���\$���E�$�����u$������  �M�l_���\$L�} ���^_���T$D����4���D$L��������A��   ����������z~�M���T$|�$R�]���D$D����$�   �$P���]����$�   Q�T$xR��$  P�Za�����P�V�H�N�P�V�H�N�P���ΉV��^������  ���؋E(�؋�Rl�D$@3�W�D$hP���ҋ�Plj�L$XQ�ˉ�$  �ҍL$dƄ$   � e���]����Dz3��}(���������D$@�#�L$d�ee���]����Dz3Ƀ}(�����L$@�   �L$T��d���E��������D�I  �D$@���/  ���&  �D$@   �M,�T$@�QR���   ��$<  Qjj���\$���E�$�ҋ�����   ��$�  P��$�   �1[����$�  Q��$   �[����$|  R��$�   �	[����$d  P��$�   ��Z����$L  Q��$�   ��Z��V��$�   R��$$  P��$�   Q�L$P��$�   R��$�   PQ�>h �����L$TƄ$    舝���L$dǄ$   �����t�����u���YX���ǋ�$�  d�    Y_^[��]�( �D$@   ������؍L$T��c���E��������Dz(�D$@��t��t�D$@   �����D$@   ��������������D$D����4���D$L��������A��   ����������z�M����$�   �$R�3Z���D$D�M ���D$|�$P�Z���L$tQ��$�   R��$  P�r^�����P�V�H�N�P�V�H�N�P���ΉV�\��������������3������3�� ����������̋D$�D$�L$��D$��� �������j�h�d�    PSVW�  3�P�D$d�    �ً|$ ����u+j@��������D$ ���|$t	���$m���3��D$��������D$$���   ���$V���҅�u*��u��t��Pj����3��L$d�    Y_^[��� �ƋL$d�    Y_^[��� ����������j�hK�d�    PQSVW�  3�P�D$d�    ��\$$3�;�t���)l����Pd����;ǉD$$��   ;�t���.h�   �������D$;ǉ|$t	����t���3��D$�������D$$P���Rm����u?�L$$;�t��Bj�Љ|$$;�u;�t��Bj����3��L$d�    Y_^[��� �ƋL$d�    Y_^[��� �ǋL$d�    Y_^[��� �V���de�  �D$t	V�U�������^� ������������V���P0j�ҋD$P����  ��^� ��U����j�h��d�    P��h  SVW�  3�P��$x  d�    ���|$P�](���D$ �D$L    u�\$L�E�    �]����D��  �E������D$ �D$ �D$ �D$ �c  �$�Ls�D$��D$�D$�
�D$�D$�u��PlV�L$0Q���ҍL$tǄ$�      �LJ���L$TƄ$�  �{Q���L$d�rQ��h��jj��$0  P�̡��h��jj��$�  Q趡���v�����<  ���  �D$@�v����l  �T$<�L$H���  j�L$0�T$H��I��� �]����Auj�L$0�I��� �]����Azj�0j �L$0�I��� �]����z'j �L$0�I��� �]����uj �L$0�pI��� �]j�L$0�`I��� �]����Auj�L$0�II��� �]����A{6j �L$0�2I��� �]������  j �L$0�I��� �]������  ����   V���҅��w  ��   +ƉD$P�Bt���Ѕ��D$$~��   Q��������D$��D$    �D$�L$��RxPQ���҅�u�D$$j �L$0�H��V�L$X���eP���j��L$0�vH��V�L$h���JP���3��9t$$�t$(��  �} �;��  �D$�D����\$��$�   ���$�	Z��3��������D$ �v  ��I �;�h  �D$P�L$X��O���D$ ���L$|��$���$��G���L$�Q�L$X�O���T$R�L$h���O����|$ �u�|$ ��  �t$P�D$\����   ��$�   Qj��$,  Rjj���\$���D$x�$�Ѕ���  �D$l����   ��$�   Pj��$�  Qjj���\$��݄$�   �$�҅��r  �|$ ��   �t$@���cT����4�L$<���$V��$   P�%P�����V����u�   �  �|$ �  �t$D���T����4����$�   �$VQ�L$X��O�����dV������   �|$ ��   ��$�   �M����$�   �M����$�   �M����$�   �M���L$H��$�   R�T$@��$�   PQR��a �T$T��$�   P�D$T��$�   QRP�a �� ��$�   Q��$�   �mO���],����z�   �:�|$ t=��$�   R��$  P��$�   �O�����!T���]4����Au�   �E�D$��D$ �t$(�����D$ �������;t$$�t$(�;����D$��tP���������E�M �    ��D$�L$tƄ$�   �'����L$,Ǆ$�  ���������D$��$x  d�    Y_^[��]�4 �I �m�m�m�m�m��V�t$W���T$���T$���$��L���D$j j V���\$���D$,�$�����_��^� �����������̃�0V��L$��K���L$��K���D$@�D$T�L$P�T$LPQR�T$T�D$P�L$,QR���\$���D$`�$�����^��0�  ����������UW�|$j ��h � @���Jz������tj j�����������tm�ESVP��������3ۅ�t?;]}:�E�<� ��tj���������t�M��R�������j �����������u��������u	^[_3�]� ��^[_]� ��������������̃�$SU3�W�ىl$�l$$�l$�l$(�l$,�-����|$4�D$(P�L$Q�������;��  3��|$ � @��;���   �T$$R�D$P��������;ŉD$ ��   �|$��   V�L$Q��� �����;���   �T$R�������D$;�|;C�C���"���3�;|$}k;�tg�L$8�D$ P�l$$������;�tG�|$ u@�L$Q�L$<�l$质���T$R�������K���S��9,�u�L$;�t	��Pj�҃�;�u��|$8^��������u_]3�[��$� �l$ ��D$ _][��$� �U����j�h��d�    P���   SVW�  3�P��$�   d�    ��}��PlW�L$XQ���ҍL$TǄ$       �C�����2  ��P4���҃��   ��Pt3ۅ��Ë�S�\$,�ҋ�����   S�Ή|$L�҅�����  ����  ��W�L$4�������Ƅ$   |
;|$<�|$8�D�D$,�D$,��$�   ����ݜ$�   �H����$�   �H����$�   �K����$�   ��J��3��L$l��$�   ��$�   �|$|��$�   �A��9}Ƅ$   �D$dt�L$T�T$\�L$P�T$L�؉D$D��L$\�T$d�\$T�L$D�T$P�D$L�D$4�L$(��RxPQ���҅���  �|$H �|$(�-  ���$    �D$4�D����\$�L$|���$�bR���|$, �D$@    ��   �D$@���L$t܌$�   �$�u@���>�\$d��$�   Pj ��$�   �ǰ   �cG���L$X��Pjj���\$����$�҅���   �>�D$|Pj ��$�   �ǰ   �#G���L$T��T$LP�jj���\$����$�Ѕ���   ��$�   Q��$�   Rj j�Ak ������   �D$@��;D$,�D$@�"����|$(��;|$H�|$(������L$lƄ$   �;����L$0Ƅ$    �j*���L$TǄ$   ���������   ��$�   d�    Y_^[��]� �L$lƄ$   ����3�9t$<Ƅ$    �D$0%tD�D$4;�t<VP�L$8�%�t$4�t$<�t$8�"�L$lƄ$   蝍���L$0Ƅ$    ��)���L$TǄ$   �����x���3���$�   d�    Y_^[��]� ��������������U����j�h�d�    P���  SVW�  3�P��$�  d�    �ى\$4��Ptj �ҋ���Ptj���҃�	����
  ��$�   �   ���AE������y�$�   �   ���&E������y�$T  �   �����	E������y�$d  �   ��I ����D������y�$�  �   ��I ����D������y�$$  �   ��I ���D������y�$  �   ��I ���D������y�$d  �   ��I ���iD������y�$  �   ��I ���ID������y�u���,  ��
�#  ��Plj �L$@Q����j�L$@Ǆ$      ��<��� �E��������Dz1j �؍L$@�<��� �T$tj�L$@�\$p�<��� ݔ$�   �\$|�ݔ$�   �T$|�T$t�\$l��Plj��$�  Q���ҋ�L$<�P�T$@�H�L$D�P��$�  �T$H����j�L$@�=<��� �E��������Dz.j �؍L$@� <��� �T$dj�L$@�\$P�<��� �T$\�\$T��T$d�T$\�T$T�\$L�L$<Ǆ$   ����諊���)�Eݔ$�   �T$|�T$t�\$l�E�T$d�T$\�T$T�\$LV�*����H������v  �����$�h�3���$�   �d$ �D�L�L$4j �~WS���\$݄�   �$�K�����ti��t'�E ���$�S�R��$8  P���gD������J����t>������|��E ���$��$�   Q��$�  R��$�   �-D�����J������  2���$�  d�    Y_^[��]�@ 3۾�����U�D�LR�{W��4t  P��4  Q�L$D��4�   P���\$݄ܐ   �$�_�����t�����   �E ���$��4�   P��$�  Q��4�   �C�����J�����a����E(���$��4�   R��$�  P��4  �ZC������I�����-����E(���$��4\  Q��$  R��4|  �&C�����I�������������H�������E ���$��$�   P��$�  Q��$�   ��B�����mI����������E(���$��$�   R��$�  P��$L  �B�����9I����������E(���$��$\  Q��$(  R��$�  �|B���J���3۾�����U�D�LR�CP�D$@��4D  Q�L$@��4�  P��4�  P��4�  P��4$  P��4�   W���\$݄ܜ   �$��������������3  �E ���$��4�   P��$X  Q����A�����oH����������E(���$��4�   R��$�  P��4  �A�����;H����������E(���$��4\  Q��$�  R��4|  �~A�����H�����Q����E0���$��4l  P��$P  Q��4�  �JA������G���������E0���$��4�  R��$�  P��4�  �A�����G����������E0���$��4,  Q��$�  R��4L  ��@�����kG����������\$8����H�S����E ���$��$�   P��$�  Q��$�   �@�����'G�����q����E(���$��$�   R��$�  P��$L  �j@������F�����=����E(���$��$\  Q��$   R��$�  �6@�����F�����	����E0���$��$l  P��$h  Q��$�  �@�����F����������E0���$��$�  R��$�  P��$  ��?�����WF����������E0���$��$,  Q��$  R��$|  �?���h���3�������D�Lj �~W��$  P���   Q�L$D���\$݄�   �$�j������4�����tV�E ���$���   P��$�  Q���   �)?�����E�����������  R��   �6?���]8�������������H���\����E ���$��$�   P��$p  Q��$�   ��>�����NE�����������$  R��$P  ��>���]8�����?  �q������D$33۾�����U�D�LR�CP�D$@��4D  W��4�  Q�L$D��4�  P��4�  P��4$  P��4�   P���\$݄ܜ   �$�������� �����4  R��4�  R����  P��$�   ����  Q����  P��$�   ����  Q��44  PW��4�  P��4�  P��4�  P��48  P�� ��0����   �E ���$��4�   R��$�  P��4�   �=�����D�����U�����4  Q��4   �=���]8�����3����E@��$�   ��$�   ��(�\$ ݄�  �\$݄��  �\$[�\$��\$� �$�o�����(��������E ���$��$�   Q��$@  R��$�   ��<�����hC�����������$  P��$P  ��<���]8����������E@�\$3��(�\$ ݄$  �\$݄$�  �\$݄$$  �\$݄$�  �$�������(���G����\$8����H��������$�  d�    Y_^[��]�@ �I �|�})��K� ���̋D$V��3�;��do�N�N�N~P��蜭�����Lf^� j�h8�d�    PQVW�  3�P�D$d�    ��t$�Lf3��|$����9~�D$�����dot�F;�tWP���po�~�~�~�L$d�    Y_^����������S�\$UVW���������GP��������o3���~6�O�<� ���D$    t� ��ȋB�ЉD$�L$Q���������;�|�_^]�   [� ���������V�������D$t	V��������^� ��V�t$��thp����k�����t��^�3�^���������������̸p�����������̋T$��|;Q}�A�I�@��� 3�� ������������VW�|$��F�NPQh�fW�������~}h�fW������_^� �V�F�Nh�fR�Vj�@PQRj j���t���_^� ���������������VW��F�N�VP�Fj�@PQR3�Wj�O ����t�F�F9F�G}��_^� �A3�9T$��R�T$R�T$R�QP�Aj�@P�ARPj j�.�����(��� �����S�\$��UV��t�L$�C����u3ۋL$��~��3�9n~<W3���L$�F�T$QSR�P�FjPj j耆���� ��t�   ����;n|�_^��]��[� �������������VW�|$W���B����~ ~�~ ~�N��X�W��6���N�VP�Fj�@PQRj j�Y �� _^� ���V��~ ~�~ ~�N��X��D$�T$PR�x6���N�VP�Fj�@PQR�AR ��^� ����������j�hh�d�    PQSVW�  3�P�D$d�    ��t$�!�  �~3ۋω\$��f��x���^�^�^9_��|�_�L$d�    Y_^[��������VW�|$��;���   SW�	�  �G�F�G�F�F�F9F �^}P������F�F��|;C�C�N�F����~"�V;Wu"�O�V�@���PQR�w
 ��[_��^� 3ۅ�~�U��I 3�9~~S3퍤$    �L$S�����N�V���ύI�ʋ��P�Q�P�Q�P�Q�P�Q�@���A��;~|���;^|�][_��^� _��^� ��������������j�h��d�    PQ�  3�P�D$d�    j$�h������D$���D$    t���>����L$d�    Y���3��L$d�    Y���������������j�h��d�    PQVW�  3�P�D$d�    ��j$��������D$���D$    t����������3����D$����tW��� ����ƋL$d�    Y_^���������������VW�|$��t5hp����z�����t%�t$��thp����b�����tW�������_�^�_2�^�������������j�h�d�    PQSVW�  3�P�D$d�    ���|$��f3ۍw�_�_�_9^�D$   |�^9^t�F;�t�SP�B���Љ^�^�^9^�\$��$t�F;�tSP����$�^�^�^���D$�����J�  �L$d�    Y_^[����������V���8����D$t	V�{�������^� ��V�t$��thx����K�����t��^�3�^���������������̸x������������VW�|$j��j���������t\�FP��������tM�NPQ��������t>���   R��������t,��   P���˿����t�NQ���������t��(V������_��^� ����̃�VW�|$��D$P�L$Q���D$    �D$    �T�����tj�|$uc�VR��������tT�FPP��華����tE���   Q���-�����t3��   R���+�����t!�|$|�FP���5�����t��(V��薶��_��^��� �����������V��W���   ���=����uj ���   PW�N�Yl�����r=���Ѕ���   �|$ ��   �L$��tA������z��݆�   �Y����z	݆�   �Y݆�   �Y����z	݆�   �Y�L$����   ݆�   �����Au݆�   �݆�   �Y����Au	݆�   �Y݆�   �Y����A��uP݆�   _�Y^� �D$��t��݆�   �X݆�   �X�D$��t݆�   �݆�   �X݆�   �X��_^� 3�9A��� �����S�\$VWS���Q���S�N�Xk������t��   ��tS�NP�	�������   �nw����_^[� ������S�\$U�l$VW��SU�O�(k������tA��   ��tSU�OP�K
������t$���   ����;����tSU���x��_^]��[� _��^][� �������j�h_�d�    PQVW�  3�P�D$d�    ��t$��  3��N�|$�dg��q���F��~�~ �~$�F(�H�~,�~0�~4�F8�H�~<�~@�~D�NP�D$� �����   �D$�u����   �~H�ƋL$d�    Y_^�������SV��W�s83�9~t�F;�t�WP�B���Љ~�~�~9{4�s(t�F;�t�WP�B���Љ~�~�~9{$�st�F;�t�WP�B���Љ~�~�~9{�st�F;�t�WP�B���Љ~�~�~�{H��   _^���   [�u�������̃�SU�ًk��VW�l$~
;k �D$t�D$ �CH��~��~	;�}9k@t3��t$U��h�gV�D$� ��������v���3���~x3�Wh�gV�����C���P��貿���|$ th�gV������K̓�Q���p����|$ t�S<�< th�gV蕼����h�&V臼��������;|$|����1���_^][��� �������j�h��d�    PQ�  3�P�D$d�    h  腽�����D$���D$    t���k����L$d�    Y���3��L$d�    Y������������SU�l$��;�t|VW�����U����  �EP�K��o���S8�R�K8�E8P�ҋC(�@�K(�U(R�ЋS�R�K�EP�ҋEH�CH�uP�{P�    󥍵�   ���   �   󥋍   _��   ^]��[� �j�h��d�    PQSVW�  3�P�D$d�    ���|$�dg�D$   �#������   �D$�Cs���OP�D$�6s���w83�9^�D$��Ht�F;�tSP����H�^�^�^9_4�w(�D$��Ht�F;�tSP����H�^�^�^9_$�w�D$��t�F;�tSP���$��^�^�^9_�w�\$��$t�F;�tSP����$�^�^�^���D$�����2�  �L$d�    Y_^[������������������j�h+�d�    PQVW�  3�P�D$d�    ��h  �A������D$���D$    t���'������3����D$����tW��������ƋL$d�    Y_^������������VW�|$��t5hx����ʇ����t%�t$��thx���貇����tW���v���_�^�_2�^�������������V��������D$t	V苼������^� ��V�t$��th�����[�����t��^�3�^���������������̸�������������V�t$��thp���������t��^�3�^���������������̸p������������V�t$��thX����ۆ����t��^�3�^���������������̸X������������V�t$��th@���蛆����t��^�3�^���������������̸@������������V�t$��th(����[�����t��^�3�^���������������̸(������������V�t$��th���������t��^�3�^���������������̸���������������������������̋D$�A� �����̋D$�A� ������V�t$W�y�    �_^� ����������̋��   �@���   ����������������́��   镼������̍��   ���������́��   �u�������̃|$ �����   � ��������������̃y �u�D$��thDhP�ն����2���� ���������̋D$hphP豶����� �����������V�t$Wj ��j��荺���O����trQ��軴������tc�GP���y�������tQ���   Q���t�������t<���   R���/�������t'���   P����������t���   Q���T�����_^� ������������VW�|$W������W�N����_��^� �hB���   �0�������������������j�hX�d�    PQV�  3�P�D$d�    ��L$�ò���~�D$    uh�   h�h�D$P�jRh�h�L$Q蓼�����L$�����P���   諺���L$�D$����花���L$d�    Y^������������VW�|$W���r�����t0݆�   �����$�۴������t݆�   �����$�������_^� ���������j�h��d�    PQV�  3�P�D$d�    ��L$�ӱ��h�   �D$h�hP�D$     跻�����L$����P���   �Ϲ���L$�D$����记���L$d�    Y^����������������VW�|$W��������t@���   P����������t+���   Q���K�������t݆�   �����$�ѳ����_^� ���������V�t$��th����������t��^�3�^���������������̸�������������j�h��d�    PQV�  3�P�D$d�    ��t$�3����N �D$    ��h荰���ƋL$d�    Y^�������������j�h��d�    PQVW�  3�P�D$d�    ��t$��h�~ ���D$   �O������D$ �C������D$�����T����L$d�    Y_^�����S�� ��5�����t�D$��thiP讲����2���[� ��[� �����������V��W�N �����|$Ph0iW�t�������V���F���h�&W�[�����_^� ���VW�|$j ��j���=�������t �FP���K�������t�� V���	�����_^� ̃�SV��^ W���N����|$�D$P�L$Q���D$    �D$    ������|$��u*��t(��V�����������tS������_^��[��� 3�_^[��� ����������V�t$��th���������t��^�3�^���������������̸�������������U����j�h�d�    P��pV�  3�P�D$xd�    ��t$@��  ����T$�T$�N�$Ǆ$�       �Ti�B"������T$�T$�N �$�*"���ƋL$xd�    Y^��]��������VW�|$��;�tPW�~�  �G�F�O�N�W�V�G�F�O�N�W�G �V��N �P�V$�H�N(�P�V,�H�N0�P�V4_��^� �������������S�A P����!&����t�D$��th�iP�*�����2���[� ��[� �������V�t$Wh�iV����������GP���ϲ��h�MV�������� W��趲��h�&V�˯����_^� ���VW�|$j ��j��譳������t �FP��軯������t�� V��詯����_^� ̃�VW�|$��D$P�L$Q���D$    �D$    �t����|$��u,��t*�VR���[�������t�� V���I���_��^��� 3�_^��� ���̸   �����������3�9D$S�\$V��W�|$��NPWS�o��Pjjj j��t������ ��t jWS�N �K��Pjjj j�t���� ��_^[� ̃�S�\$ VWS���~{���wV�D$P��辬�����P�V�H�N�P�V�H�N�P�V�w V�D$P��茬�����P�V�H�N�P�V�H�N�P_�V^�   [��� ������������SU��V3�W�]�}�    �hY󥍍�   ���   ���   ���   ��������   ����_^���   ][����h�7���   ��������������������U������   �} SVW��u"�E� F�P�P��E��i�P�P��L$�����L$@�E����~@W�^(�D$,SP�c'����h(�h�h��h�=�L$8QWS�VR�L$`����3�9��   ��   3����    ���   �P�L$�^"���M�A�D$��������z�Q�A�D$ ��������z�Q�M��D$��������Au�����A������z���Y����Q����Au�Y��؃���;��   �o���_^�   [��]� ̋��L$��|;��   }����   �T$R���� ��������j�hK�d�    PQ�  3�P�D$d�    j(�X������D$���D$    t���N����L$d�    Y���3��L$d�    Y���������������j�h{�d�    PQVW�  3�P�D$d�    ��j(�������D$���D$    t����������3����D$����t;�tW����{���� W�N �@����ƋL$d�    Y_^���������������VW�|$��tEh�����Zy����t5�t$��t-h�����By����t;�tW���r{���� W�N �֮��_�^�_2�^�������������V�������D$t	V��������^� ��j�h��d�    PQ�  3�P�D$d�    j8�ث�����D$���D$    t�������L$d�    Y���3��L$d�    Y���������������j�h��d�    PQVW�  3�P�D$d�    ��j8�d������D$���D$    t���������3����D$����tW��� ����ƋL$d�    Y_^���������������VW�|$��t5h������w����t%�t$��th������w����tW�������_�^�_2�^�������������V���Ti�R�  �D$t	V襬������^� ������������SUV�鍵�   3�9^Wt�F;�t�SP�B���Љ^�^�^���   �W������   �L����]�}�    �hY�_^���   ][����������������j�h=�d�    PQVW�  3�P�D$d�    ��t$�2�  3��N�|$�j����ǆ�   lI���   ���   ���   ���   �D$蒥�����   �D$肥�����D$�6����ƋL$d�    Y_^�����j�h��d�    PQSVW�  3�P�D$d�    ���|$�j�D$   �������   �D$�3������   �D$�#������   3�9^�D$�lIt�F;�tSP���xI�^�^�^�O�\$��_�����D$�����v�  �L$d�    Y_^[������SU�l$��;�taVW�������F���U����  �E���   �R�C�u�{�    󥍋�   ���   P�ҍ��   P���   �������   _���   ^]��[� ������������U������VW�������}�D$P�L$Q���D$    �D$    �ڪ���ȅ���   �|$��   �T$R���ؓ���ȅ���   �D$P�c������NQ�ωF�����ȅ�t`���   R��譜���ȅ�tK���   P���x����ȅ�t6���   Q���c����ȅ�t!�T$R���`����ȅ�t�|$ �����   �F���xj��������{a�F��������AtS�F ��������AtE3�9��   ~/���   ���������At(�G��������At����;��   |׋���_^��]� _��3�^��]� ��������V��������j��^�����������������j�%��������V���x�����j��^�����������������j����������V���H�����ݖ�   �tkݞ�   ��^��tk����������VW�|$W��������ȅ�t&���   P��螒���ȅ�t���   Q��艒������ܖ�   ����t8�xjܖ�   ����{#��ܞ�   ����tܞ�   ����{_��^� ����_3�^� ������j�h��d�    PQV�  3�P�D$d�    ��t$�c������   �D$    ��k�J������ݞ�   ǆ�   �  �ƋL$d�    Y^����j�h�d�    PQVW�  3�P�D$d�    ��t$��k���   ���D$   ��������D$ �������D$�����a����L$d�    Y_^������������������VW�|$��;�t2���   P���   �B������   ���   ݇�   Wݞ�   �������_��^� �����������VW�|$W���"����ȅ�t;���   P���.����ȅ�t&���   Q���)����ȅ�t���   R��褐����݆�   _��^�xj����Au3�� ��� V��������dl��^����������������dl�U��������j�h;�d�    PQV�  3�P�D$d�    h�   褣�������t$3�;��D$t���j�����j�ƋL$d�    Y^����j�hk�d�    PQVW�  3�P�D$d�    ��h�   �A��������t$���D$    t��������j�3����D$����t;�tW���C����ƋL$d�    Y_^������������������VW�|$��t9hp����o����t)�t$��t!hp����o����t;�tW�������_�^�_2�^���������j�h��d�    PQV�  3�P�D$d�    h�   �d��������t$3�;��D$t���*�����j�ƋL$d�    Y^����j�h��d�    PQVW�  3�P�D$d�    ��h�   ���������t$���D$    t���������j�3����D$����t;�tW�������ƋL$d�    Y_^������������������VW�|$��t9hX����zn����t)�t$��t!hX����bn����t;�tW������_�^�_2�^���������j�h��d�    PQV�  3�P�D$d�    h�   �$��������t$3�;��D$t���������ݖ�   �tkݞ�   �ƋL$d�    Y^������j�h+�d�    PQVW�  3�P�D$d�    ��h�   豠�������t$���D$    t���u�����ݖ�   �tkݞ�   �3����D$����t$;�t W������݇�   ݞ�   ݇�   ݞ�   �ƋL$d�    Y_^������������VW�|$��tQh@����
m����tA�t$��t9h@�����l����t);�t W���2���݇�   ݞ�   ݇�   ݞ�   _�^�_2�^�j�h[�d�    PQ�  3�P�D$d�    h�   襟�����D$���D$    t��������L$d�    Y���3��L$d�    Y������������j�h��d�    PQVW�  3�P�D$d�    ��h�   �1������D$���D$    t���g������3����D$����t6;�t2���   P���   菡�����   ���   ݇�   Wݞ�   �������ƋL$d�    Y_^��������������VW�|$��t5h(����k����t%�t$��th(����rk����tW������_�^�_2�^�������������j�h��d�    PQV�  3�P�D$d�    h�   �4��������t$3�;��D$t��������dl�ƋL$d�    Y^����j�h��d�    PQVW�  3�P�D$d�    ��h�   �ѝ�������t$���D$    t�������dl�3����D$����t;�tW��������ƋL$d�    Y_^������������������VW�|$��t9h����Jj����t)�t$��t!h����2j����t;�tW���r���_�^�_2�^���������V�������D$t	V��������^� ��V����j�r����D$t	V��������^� ������������V����j�B����D$t	V赞������^� ������������V���tk�����D$t	V腞������^� ������������V���(����D$t	V�[�������^� ��V���dl������D$t	V�5�������^� ������������V�t$��thЉ����h����t��^�3�^���������������̸Љ�����������V�t$��th�����h����t��^�3�^���������������̸�������������V���ط  3��F�F�FL�FP�F�F�F�F�F �F$�F(�F,�F0�F4�F8�F<�F@�FD�FH��n��^���̸   ����������̃yP u3�� �y4 t��y8 t�y< t�V�q��|�A��|�Q��}3�^� S�Y;�}[3�^� W�y ;�|�A$;�|�q��~�Q��t��t_[3�^� ��U�nu��QL��~������;�|Q�A@�qH3�;AD�   ��+�;t�@}�؋º   �;t�@}	�ظ   ��   �|�@;�|�T��t�@��;�}	]_[3�^� �D���3�9D�@]��_[^��� ����������SV���P0j�ҋFP3�;�t9^L~P�o������^P�F4;�t9^(~P�W������^4�F8;�t9^,~P�?������^8�F<;�t9^0~P�'������^<�^L�^(�^,�^0�^@�^D�^H�^�^�^�^�^^[����������̀y t�A��~��ËA�����������̋AP��t$�Q@�T$V�qD�t$�IH�L$�э�^� 3�� �APS2ۅ���   �Q@�T$V�qD�t$֋qH�t$֍Ѕ�^��   8YtR�A��������D{q�A���4D$�����y~�B������X�y~��[�J�X�� ��[�X�� ��D$��y��~�B����X�y~���B�X�[� �؊�[� ������������VW�|$����~A�NL;�}:�FP��t��t/��    QP�Ĳ�������    R�R������FP���#ǉFL�~P _��^� �������VW�|$2�����wWS�\$��~M�L�(;�}=�D�4��t��t1��    QP�V��������    R�������D�4���#ÉD�(�|�4 ��[_^� �����V��F�P�N�ҋF8�P�N8�ҋFx�P�Nx�ҋ��   �P���   �ҋ��  �P���  �ҋ�^�d����V��N����Wth��t8��t �D$3���tQh,oP�ҕ������_^� ���  ���  _^�@���Vx�|$�B�NxW�Ѕ�tԋ��   �B���   W��_^� �V�|$�B�NW�Ѕ�t��V8�B�N8W��_^� �����V�t$W���GPhhoV�I���hToV�>�������贔���G��t`��t1��un��  Q���d������  �B���  V�Ћ�軔��_^� �Wx�B�OxV�Ћ��   �B���   V�Ћ�葔��_^� �W�B�OV�ЋW8�B�O8V�Ћ��m���_^� �������̸   �����������V��F8�P0W�|$�N8W�ҋ��   �P0���   W�ҋ��  �P0���  W��_^� ��̋Q3���t,��t��u-���  �P4���  �⋁�   �P4���   ��A8�P4��8����������������̋Q3���t$��t��u$���  ��@8�����   ��R8���8��@8��� ����̋Q2���t0��t��u8���  ��T$�@<�����   ��D$    �R<���8��D$    �@<��� ̋Q3���t$��t��u$���  ��@D�����   ��RD���8��@D��� ����̋Q3���t,��t��u-���  �PT���  �⋁�   �PT���   ��A8�PT��8����������������̋A��t)��t��t3�� ���  ��@X�����   ��RX��A8�@X��8�����̋Q2���t%�I��~V�t$��t��~VjPQR�HE�����^� ��������������̋Q2���t%�I��~V�t$��t��~VjPQR��D�����^� ���������������j�h!�d�    PQ�  3�P�D$d�    �L$�L$���D$    t��� �L$d�    Y��� ����j�hK�d�    PQ�  3�P�D$d�    jT��������D$���D$    t���>����L$d�    Y���3��L$d�    Y���������������U����  3ŉE�SVW�}j j��h � @����0�����  �CP���e������E���   �KQ���N������E���   �SR���8������E���   �CP���"������E���   �KQ���������E���   �SR����������E���   �C P����������E�tw�K$Q���Ύ�����E�te�S4�C�KRPQ�FG ��P��軎�����E�tB�S8�C �KRPQ�#G ��P��蘎�����E�t�S<�C$�KRPQ� G ��P���u����E��{ t�s���u���S�U���    �=� ���ĉE�~�5������������x�}�{ �E�    ��   �}� ��   �{  �E�    ~d�}� t^3�9s$~I�}� tC�CP��t"�KH�SD���U�}ʋS@�U�ʍȅ�u�E�P�E�P��赍����;s$�E�|��E��;C �E�|��E���;C�E��s������c�����u���e�_^[�M�3��� ��]� �E���j�hx�d�    PQV�  3�P�D$d�    ��t$��n�D$    ��������D$����趬  �L$d�    Y^�������̃�0U�l$<��VW�|$@��t�������u	3����F���L$H����   ����$�ύ������   �L$������~ �D$D    ��   S3�9^ �~   3�9~$~o�L$H�D$PWSQ���6����L$L�T$R�D$,P�S�����L$�P�T$�H�L$�P�T$�H�L$ �P�L$DU�D$P�T$,��L����t�   ��;~$|���;^ |��D$H��;F�D$H�c���[_��^��]��0� UW��膰  ��t�   _��^��]��0� ��������������̃�SUVW���\���N���FPQ��L� D �V ��FRP�D �N$�VQR�D$,� D ���~ �D$t�F��~����F�^ �N$�V������L$L$͍�_^][����������������QUV��L$W�FPjQ��  �VRjP��  �NQjP��  �~WjP��  ����0����   �~  ��   �V$����   �~@ ��   �~D ��   �~H ��   �~P ��   S����������D$�3ۅ�~i3�9F �D$~S��I �~P��t�ND�ȋF@��ȍ<��3�;�}�L$WQU���  �VH�<׋V$��;ڋ�|�D$��;F �D$|���;^�~|�[�F4��VPQR�B �����PU��  �N �V�����F8PQR�pB �����PW��  �N���F$PQ�QB �V<��R�PW�`�  �� _^]Y� �����́�   �  3ĉ�$�   SUV��$�   W��F$�N �VP�FQ�NR�VP�F�~Q�NRPQh�oh�oS������,3퍛    ��w��G�RP�A ���3�PUh�.S�ۊ���O��G��QRP��膕��������|��~ ��<u��<�N �N�N$PQh�<S蓊�����~P uhx<S�������   h�   �T$j R��� 3��9n��   3�9~~r�����~h�&S�=�����WU�D$h�oP�D$  ��� �FP����t�ND�V@����ʍ��3��VH�L$Q�NP�F$R�VPQR���w�����;~|��F��;�}h�&S�ʉ������;n�c�����$�   _^][3��� �Ą   � SV�������\$���L$�D$��  ����  ����  9\$ W��  �|$(;���  �T$,;���  �L$��}$h�ph�ph#  ho������_^2�[�  �D$<t��th\ph�ph)  �΄����F����FH�FD�ǉ^�\$�^�\$ �^�\$$�F@�ÉNP�Ή^�~ �V$�����N�VQR�~? ��Pj ��������F �NPQ�d? ��Pj��������V$�FRP�J? ��Pj��������N4�V�F���$QRP�TM ��N8�\$�V �F��QRP�:M ��N<�\$�V$��QR�FP� M ��N4�\$��V�F�\$��QRP��E ��N8�\$��V �F�\$��QRP�E ��N<�\$��V$�F�\$��QRP�E ��B��j ����_��^��[�  h0ph�ph  �^����|$ u,�|$ u%��u!��u��u9L$ u9L$$u9L$(u^�[�  hph�ph  ho�7�����^2�[�  �������������QSV��~P ty�   9F|o9F |j9F$|e�~@ ~_�~D ~Y�~H ~S�L$U�l$��D$    W�	��$    ���T$;V��   3���t};~ }x�FP��t<�VD�^@���\$Ӎ��)h�ph�ph�  ho2�������^��[Y� 3�3҅ɋL$��R�VHUQ�NP�F$R�VPQR�nL���   �� ���u��D$���c���_]^��[Y� �������̃�V��~ ��  ��P4U�ҋ�F����  �V ����  �N$����  ����  9n@SW��   9nD~9nH~z���D$    ~[��3�9V ~@3�9F$~1�NP��t�~H�^D������^@�\$����3Ƀ���;F$|σ�;V |��D$��;F�D$|���_�F�~ []��^��Í]�����������W�\$ 谠�������~ ��    �|$ �D$�D$    ��   3�9n �l$~c3�9^$~L�FP��t!�NH�VD���Ջl$ʋV@�T$ʍ��3��L$QPW�r� ��|$ �������;^$|���;n �l$|��\$�D$��;F�D$|��|$ �V$���V �VR���F�^����F$���F �F�NP���PWQ��� W�	����F$�V �Ã���_�^H�FD�V@[�~ ]��^�����VW���G�P�O�ҋ��G8�P�O8���   �ҍOx���P�ҍ��   ���P�ҍ��  ���P�ҋ�  �����_�^��QV�t$Wjj��h � @���w#����u_3�^Y� �GSP���߁���؄���  U3�Ujh � @���C#���؄��  �G��t!��t��u'��  Q���I�������Ox��O��B V�Ѕ��Ë��i�����u2��4  ���,  Ujh � @����"���؄��  �G��t��t��u ���  ����   ��O8��B V�Ѕ��Ë�������u2���   ����   V���  �E9���؄���   Ujh � @���\"���؄���   ��  P�ΉD$�����9l$��~,�l$�d$ ��t ��  L$V蜵 �D$P��;l$��|܋��u�����u2��C��t?݇  �����$�����؄�t&��   Q��葪���؄�t��!  R���|�����]���"�����u2���[_^Y� �̃�0UVW��������t$@�D$8P�L$4Q3�h � @�Ή|$<�|$D�_������k  �|$0Sth@rh,rj%�  �T$,R�Ή|$0�|$ �|$�|$(�|$�|$�|$$�|$,�n���؄���  �D$,���='  ��  �L$(Q���zn���؄���  �D$(;�t��thrh,rj>�  �T$R���Fn���؄���  �D$���='  �`  �L$Q���n���؄��s  �T$�����'  �)  �D$$P����m���؄��J  �L$$�����'  ��  �T$R����m���؄��!  �D$;D$��  =�� ��  �D$P���m���؄���  �D$;D$��  =�� �x  �L$ Q���nm���؄���  �D$ �L$$;��D  =�� �9  �T$�|$(P�D$R�T$$PQ�L$(Q�L$@��RPQ���>����؄��s  �U4�E�MRPQ�6 ��P���m���؄�t@�U8�E �MRPQ�q6 ��P����l���؄�t�U<�E$�MRPQ�O6 ��P����l���؀} t�E���D$8��U�T$89|$�|$0��   �L$�D$ ��3�����   ��~O����tI3���~8��    ��t*�D$0VWP��������L$8PQ�L$L�Ol���؋D$ ��;�|ҋL$�t$D��;�|��T$0��;T$�T$0|��oh�qh,rjz�Rh�qh,rjp�Dh�qh,rjf�6hlqh,rj\�(hHqh,rjR�h$qh,rjH�h qh,rj4ho�V�����2ۋ�������u[_^��]��0� ��[_^]��0� _^��]��0� V�������D$t	V�k�������^� �̃�SUVW�|$ ��;��  W�ś  �G$�O �WP�GQ�OR�WP�GQ�ORPQ���-�������  �C��|1�K;�|*�{4 t$�4 tQP�s4 �W4���P�C4RP�/� ���C��|1�K ;�|*�{8 t$�8 tQP�:4 �O8�S8���PQR��� ���C��|1�K$;�|*�{< t$�< tQP�4 �K<���P�G<PQ�� ���{P �3  �GP���D$ �$  �S@���  �{D �  �sH���  ������;W@�,�    �l$u9�CD;GDu1;wHu,�S$�S �S�D$ ��RP�CPP�@� ��_^]��[��� �{ �KP�L$ �D$    ��   ���    �{  �D$    ~b�C$3���~I�GP��t#�WH�OD���L$�l$ыO@�L$э��3��T$ UPR��� �C$l$,����;�|��L$��;K �L$|��D$��;C�D$|�_^]��[��� �������_^]��[��� ���SV��~ W~�~  ~�~$ t�|$���|$�����$2���z������   ��~ u2�W`����Dz�Wh����Dz�_p����D{���7���������,������U3��ta�;n}[3���tN��I ;~ }D�FP��t�ND�V@����ʍ��3��L$�VHQ�NP�F$R�VPQR�s �؃�����u�����u�]_^��[� _^��[� �������������SUVW�|$����}S3�9n�
  �~��x"�������    �N��� ����P;�}�N��PUQ����_�n�n�n^][� �F;�}k�N��PWQ����3�;ŉF��   �V��+ʍ�����Q���UR迻 �F��;�}������+�F�P���������P��u�~_^][� ~T���;�|%��+������荛    �N��&� ��P��u�9~~�~��F�RWP�Ή~��3�;ŉFu�n�n_^][� ���������������j�h��d�    PQVW�  3�P�D$d�    ��jT�z�����D$���D$    t����������3����D$����tW��� ����ƋL$d�    Y_^���������������VW�|$��t5hЉ���:G����t%�t$��thЉ���"G����tW�������_�^�_2�^�������������UW��3�9o�|ot7V�w��xS�����O��� ����P;�}�[�O��PUQ���҉o^�o�o_]����������������U�l$V��;�tX�ES3�;��^[��^]� 9F}P�d���9^t�E;ÉF~�W3����E�N�P���� ����P;^|�_[��^]� ��^]� ����̋D$9A}	�D$����� �����������UW��3�9ot<V�w��x!S������I �O���� ����P;�}�[�O��PUQ���҉o^�o�o_]�V�������D$t	V�z������^� ��SU�l$VWU��� �  �E�MQ�K�C�N%���U8R�K8�B%���Eh�Ch�Ml�Kl�Up�Sp�Et�MxQ�Kx�Ct��������   R���   ��������   ���   ���   ���   ��   ��   ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �    ���  �R���  �g������  P���  ��,����  Q��  �����݅  ݛ  ��   _��   ��!  ^��!  ]��[� ������VW�|$��t5h�����JD����t%�t$��th�����2D����tW������_�^�_2�^�������������j�h8�d�    PQSV�  3�P�D$d�    ��t$�2�  3ۍN�\$��r�^�k ���N8�D$�^ ���Nh�D$������Nx�D$��������   �D$�����h@h`�jj���   P�D$,�
� ����$��  �D$ �]n�����  ��������  �D$�b*����ǆ  |o��  ��  ��  ݞ  ��   ��!  �ƋL$d�    Y^[�����������������j�h��d�    PQV�  3�P�D$d�    ��t$��r��  �D$   �������  �D$�*�����  �D$�?���h@jj���   P�D$$�� ���   �D$�%!���Nx�D$�!���Nh�D$�;,���N8�D$�^M���N�D$ �QM�����D$�����ґ  �L$d�    Y^����V��  �F    �{p���N�3 ���N8�+ ���Nh�c����Nx�[�����   �P�����   �E�����  �:������  �������  ������  ������ݞ  Ɔ    Ɔ!   ^��V��F�V����;�uJ��   v��|��� ;�}�������   ��;�}8P���'����N����F���N^�N�+� �F����V��R�����N����F���N^����j�h�d�    PQ�  3�P�D$d�    h(  ��s�����D$���D$    t�������L$d�    Y���3��L$d�    Y������������j�h;�d�    PQVW�  3�P�D$d�    ��h(  �as�����D$���D$    t���'������3����D$����tW���}����ƋL$d�    Y_^������������V�������D$t	V��t������^� �̃�DSVW��������|$T3��D$�D$�D$P�L$Qh � @�������؄��H  �D$��UuQ���  �B$���  W�F   �Ѕ��Ä��
  W���  �	(���؄���  ��  V���q_������  ����  �nU���6^���؄���  �L$Q�T$\3�Rh � @�ωD$d�D$�|����؄���  �|$X�Ä��  �E ����   ��t����   ��  P����^������   �Vx�B$�nxW���Ѕ��Ä���   �U �Rlj �D$(P���ҋ���   �P���   �H��   �P�L$$��  �[(���E �Plj�L$8Q���ҋ��  �P��  �H��  �P��  �L$4�A�F�P$�nW���҅��Ä�t/�E �Ph�L$DQ���ҋ�Nh�P�Vl�H�Np�P�Vt�L$D��'�����d������|  ���v  �D$P�L$\Q3�h � @�ωl$d�l$�$����؄��L  �|$Xu-�F��t��t��u���  ����   ��N8��B$W�Ћ�����W���  �&���؄���   �L$Q�T$\Rh � @�ωl$d�l$諦���؄���   �|$X�l$�Ä�t"�D$P���\���؄�t�L$Q��  ������|$ ~7�D$    ��t+��  �a�����  L$W�� �D$P��;l$��|ы��:�����tV��tT�|$ |@��  R���-\���؄�t9��   P����i���؄�t%��!  V����i���؄�t�2ۋ�������u2�]_^��[��D� �V�t$��th�����;<����t��^�3�^���������������̸�������������j�hs�d�    PQV�  3�P�D$d�    ��t$�3�  �N�D$    �ds�]�����8  �D$�]�����^�ƋL$d�    Y^��������j�h��d�    PQV�  3�P�D$d�    ��t$�ds��8  �D$   �F���N�D$ ��������D$������  �L$d�    Y^����̋�8  �P��8  ����������������́�8  ��@�����VW�|$��W�N�o�����8  �P��8  W��_^� ��������VW����;������8  �P��8  ��`  ��_�^����������V�t$Wjj��h � @�������u_3�^� Sj jh � @�������؄�tpV�O�M����Ί��D�����u2��V��tRj jh � @������؄�t<��8  �P ��8  V�҅�����������u2����t�G�����$�k���؋��ߔ����u2���[_^� ����UV��W�^�F�~�ωD$������8  �������t$ 3��D$�D$�D$P�L$Qh � @��������u_^3�]��� �|$S�Ä���   3��T$$�D$�D$$R�D$Ph � @��������؄�t{V�������Ί�躖����u2��b��t^�L$$Q�T$3�Rh � @�ΉD$0�D$�~����؄�t8�E �P$V���҅������q�����u2����t�|$|�D$P���bX���؋��I�����u2���[_^]��� �����̸ �  ����������̋�8  �P4��8  ����������������́�8  ��@8����́�8  ��@<����́�8  ��@D�����j�h��d�    PQ�  3�P�D$d�    hh  �5k�����D$���D$    t��������L$d�    Y���3��L$d�    Y������������V���8����D$t	V��l������^� ��VW�|$W���B�  �G�G�^P�N�������8  W��8  �^��_��^� �������VW�|$��t5h�����j7����t%�t$��th�����R7����tW������_�^�_2�^�������������j�h��d�    PQVW�  3�P�D$d�    ��hh  �j�����D$���D$    t����������3����D$����t,W���]�  �G�G�^P�N������8  W��8  �y���ƋL$d�    Y_^��������V�t$��th�����{6����t��^�3�^���������������̸�������������j�h>�d�    PQSVW�  3�P�D$d�    ��t$�T���~���D$    �t��[ �^8���D$�
������D$������N ���������FH   ����^@�L$d�    Y_^[����j�h~�d�    PQSUVW�  3�P�D$d�    �ى\$�pS���t$(�k�   ���t�D$     �s8���D$ �s������D$ �CH   ��[ ��;������u������\$�����$�*����ËL$d�    Y_^][��� ��j�h��d�    PQV�  3�P�D$d�    ��t$�t�N8�D$   �����N�D$ ������D$������R���L$d�    Y^����������R����H��������V��L$�FPj0Q�-�  �V8RjP�!�  ��HVjP��  ��$^� ��������������SU�l$��;�t5VWU�`���u�{�   �E8�C8�M<�K<�U@�S@�ED�CD�MH_�KH^]��[� �������̋AH������������̋T$3�9D$V����L$PQR�N�!���P�FHjjj P�+���� ��^� �������VW�|$W���R2�����{R��W�N�\ _��^� ���������̃�UW�|$3�������   S�\$��w|;�txV�uW���P���� S�\$���B���W�ΉD$ �6����L$�S����&����D$�u �W������� S�\$������W�΋�������E S���������D$��   ^[_]��� ����������̃�VW���w8j ��������\$j��������\$����Au"�O�Y ��$����Au�_��^��� 2�_��^��� ������SVW���w8j���������$j �������t$���$huV��c�������qc��h�tV��c�����_S���f��h�tV��c������ W���f��h�&V�c�������ZX ���$h�tV�c�������Oc��_^[� ���������VW�|$j ��j���mg������t2�FP���˅������t �N8Q���Ɇ������t�VHR���wa����_^� ��������������̃�VW�|$��D$P�L$Q���D$    �D$    �g������t9�|$u2�VR���Q������t �F8P���R������t��HV����O����_^��� ������������Q�D$�Q8��Q<�P�Q@�ID�P�$    �HY� ����������D$V�D$��������z$�����\$�N8�$�������aO���   ^� ��3���^� ��������������VW�|$�G�����wO9~HS���   �O���   ;�uI�F�5��������D��{�V�F ��������D{���^0[_�NH^� _2�^� ����[_�NH^� 9NHuU�F�5��������D��{�F������Dz�V�F������D{ �F0��������Dz���^[_�FH   ^� �����FH   ��[_^� ����VW�q8j �������|$j��������_������_��^� ̋�Pj ��� ����SV���PWj �ҋ|$����tB��t>�D$���~H�$Wu������_^[� �����X ��u����$��W�X ��_^[� ��SVW�D$P��3��`���|$(P��� ������\$,����Az$�L$Q���a��P���ߣ�����\$,����A�C{��_^[��� ���̃�SUV��n�F�N�V�^�l$ �n W�~�n�n$�n�n(�n�n,�n�n0�n�n4�F �D$$�N$�V(�~,�^0�N8�n�F4���������L��_^]�   [��������������U������tSVW��3ۍw8S�������\$Hj�������\$H����A�}  j��������]����Dz���.j ��������mj���\$D�����j �\$L�������l$H�|$@���D$X�$�OP�1T �D$P�u��D$X�^�Hu�D$`�^�}��   �]ۍGP�L$l�QۍO ��~���j�O8�T����\$Hj �O8�F����l$H�D$h�   ����D$p���^9GHu	�|$x�^��؋M��Q����D$@   |Z�Q����T$H��   �T$@�T$H���V9GHu�V���V9GHu�V���V9GHu�V���V9GHu�V��u��T$@;�+ʃ����V9GHu�V��u��ظ   _^[��]� _^��[��]� ̋D$�T$�A�D$�Q�T$�A�D$�Q�T$�A�Q��J���   � ��������̋D$�T$�A �D$�Q$�T$�A(�D$�Q,�T$�A0�Q4�J���   � ���������U������4SV�uW��3�3ۃHj��jS�΃�P�T	������  �_8j ���D$   �����\$j�������T$�]�D$��tj��������   ��j �����r����\$ j���e����D$�D$ ������z�����D$������z��������������zo�����T$���T$��������zd�N��V�Ƀ��Z�D$0���$P�*\��Pj �������D$���L$0�$Q���
\��Pj���`����D$_^[��]� �����D$    ���3�����AuU�V����F�Ƀ��X�L$0�$Q���[��PS�������D$���T$0�$R���[��Pj���������_^[��]� �F���؍W��R�j �N���Y��������� Wj������_^��[��]� ������������̃�0SVW�|$@���3���������   ���H��S����������D$�$P���[��j����������L$,�$Q����Z���T$$R�L$�Y�����$����Aup�D$�L$�T$�F�D$�N�L$�V�T$ �F�D$$�F �D$0�N�L$(�N$�L$4�V�T$,�V(�T$8�F,�N0�V4��F8�O�N<�W�V@�G�FD�   ����G��_^��[��0� ����������U����j�h�d�    P��(  SVW�  3�P��$8  d�    �ً�Ph��$�   Q���ҋ�Ǆ$@      �y����\$T�����$�   ��$@  �_����$�   �{P����N �W�G��T$`�W�D$d�G�L$\�O�T$l�S$�D$p�C(�L$h�K �T$x�S0�D$|�C4�L$t�K,��$�   ��Rh��$�   ��$�   ��$�   P����j ��Ǆ$D     ������ ��$�   ݜ$�   ��$@  �����Ph�L$DQ����j��Ǆ$D     ����� �L$Dݜ$�   ��$@  �u����L$DQ�D$C �ˋPh��j��Ǆ$D     �~����uj�ΉD$D�~����D$@��D$>����At�D$> �L$DǄ$@  ��������|$> ��   ��Rh�D$DP����j��Ǆ$D     �����D$@��$�   Pj�������L$D�!����$�   �t$`�$R������P�L$x�G����L$DǄ$@  �������j�������ݜ$�   �D$?��Ph�L$DQ����j ��Ǆ$D     ����j �ΉD$D�����D$@��D$>����{�D$> �L$DǄ$@  �����$���|$> ��   ��Rh�D$DP����j ��Ǆ$D     �'����D$@��$�   Pj ���"����L$D�!����$�   �t$`�$R�������P�L$`�X����L$DǄ$@  �������j �������ݜ$�   �D$?��|$? tS�D$tP�L$`Q��$�   �����   󥍌$�   �[���݄$�   �Bl�����\$݄$�   �$�Ћ��#D���D$?��$8  d�    Y_^[��]� �������j�hK�d�    PQ�  3�P�D$d�    jP�X�����D$���D$    t�������L$d�    Y���3��L$d�    Y���������������j�h{�d�    PQVW�  3�P�D$d�    ��jP�W�����D$���D$    t���������3����D$����tW��� ����ƋL$d�    Y_^���������������VW�|$��t5h�����$����t%�t$��th�����$����tW������_�^�_2�^�������������V��������D$t	V��X������^� ��U����j�h��d�    P���   SVW�  3�P��$�   d�    ���Ej�^8�����$3���������   �FHW�ˉD$4莾��ݜ$�   j���~���ݜ$�   �L$4�.I �L$d��$   �I �E�N�V�F�~�L$4�O�T$8�W�D$<�G�L$@�����$Ƅ$  �T$L�D$P�i�������$�   �$Q���I ��L$L�P�T$P�x�|$T�X�\$X�X�\$\�@�T$h�T$X�L$d�N$�D$`�T$p�V(�D$x�F ��$�   �N0�D$|�F,��$�   �V4��$�   �L$4�|$l�\$t��$�   ��$�   �H ��$����D��   �L$d�H ��$����D{k�}�7��th�����"����t�t$,��D$,    �t$,�E���th������!����u3ۃ? t_��u[h�uh�uhN  hhu�n������L$dƄ$    ����L$4Ǆ$   �������3���$�   d�    Y_^[��]� �M�9 t��uh,uh�uhS  뗅�u5jP�dT�����D$,��Ƅ$   t	��������3�Ƅ$   �D$,�����u7jP�+T������$�   ��Ƅ$   t	�������3��UƄ$   �؉����?���E�~���   �\$݄$�   �t$D��$�t$<�N8�����D$0�ˉFH�?��݄$�   ���\$�{�E�   �t$t�$�K8�~����L$0�KH�L$d�   Ƅ$    �Q
���L$4Ǆ$   �����=
���ǋ�$�   d�    Y_^[��]� ��̃�SUV�t$3�3�;�W�L$t9n|�n�|$ ;�t9o|�o��PU�҅��	  ;��   tr�F;�}M9^~�^�N��PSQ����;ŉFt*�V;�}��+ʍI���Q�R��UP�� ���^��n�n�L$��Q���ծ���T$�� R���Ʈ��;���   �G;�}G9_~�_�O��PSQ����;ŉGt$�O;�}��+����R��UP�~� ���_��o�o�t$��8U���A����\$�L$Q�����j���(����\$�T$R������_^]��[��� �����������̸�������������j�h�d�    PQV�  3�P�D$d�    ��t$�s<��3��N�D$�v�F�F艹���N �D$�|����ƋL$d�    Y^������������j�h>�d�    P��UVW�  3�P�D$$d�    ��t$��;���D$4�~���D$,    �v�F�F �����n ���D$,������N���D$,tB��Rh�D$P�ҋ�M �P�U�H�M�P�U���P�W�H�O�P�L$�W����ƋL$$d�    Y_^]�� � ���������;����(��������V��~ t�N��T$�@R����D$�NQjP���  �VRjP��  �� VjP�ި  ��$^� �������VW�|$��;�tDW��H���G�F�O�N�W�V�G�F�O�N�W�G �V��N �P�V$�H�N(�P�V,_��^� ���������j�hs�d�    PQV�  3�P�D$d�    ��t$�v�N �D$   �F    �k���N�D$ �^�����D$�����:���L$d�    Y^�����������������V��~ u�F P�N�{�����t.�D$���N �$蕷���~ t������N�$�=���^� �D$^� ̃��D$V���\$�~ u�F P�N� �����t1�D$���N�$�:����~ t������N �$����^��� �D$^��� j�h��d�    P��V�  3�P�D$$d�    ��D$8���D$    u.�N�D$4��V�P�N�H�V�P�L$$d�    Y^��(� �N �V$�L$�N(�T$�V,�L$�T$ P�L$�D$0   ����3�8F�L$��P����� �����$�����\$3�8N��Q�L$����� �����$�x����t$4���\$���D$�$�����L$�D$   �D$, �y���ƋL$$d�    Y^��(� ���̊A�������������j�h��d�    P��SV�  3�P�D$d�    ���D$$    �9���L$,�c����؄�t}�N��tZ��@h�T$R�ЍL$,Q�L$�D$(�����L$�.����؄�t�T$�D$�L$�V�T$�F�N�V�L$�D$$ �����D$,�L$0�T$4�F�D$8�N�V�F�L$,�D$$��������ËL$d�    Y^[��� ���������Q�D$�Q��Q�P�Q�I�P�$    �HY� ���������VW���O3���t[;�tW��Pd�ҋ���tJ����   �OQ���Ҁ t����   ���ҋW �G ���̉�P�Q�P�@�Q�A����7����_^������j�h�d�    P��SUVW�  3�P�D$(d�    ��l$8�D$    �~ t5�N��PU�ҋ؅�tZ�~��躴����u3ۅ�tFhtwU�%J�����63��2�N��@h�T$R��j W���D$8    �D$   蓶�����D$8t�D$8 �D$�D$0����t	�L$�����|$8 t,3���th(wU�I�����ƋL$(d�    Y_^][�� � ��t�N ������u3���t�h�v�������������V��W�~j���в�����$j ��������F�L$���$Ph�wQ�8I����_^� �y t
�I��@8��3�� �����������Q�D$�Q ��Q$�P�Q(�I,�P�$    �HY� ����������D$V�\$��3�����Au*����5���D$���\$�N �D$�$������   ^� ��^� ������������j�hH�d�    PSVW�  3�P�D$d�    ��>j�L$$�D$    趱��j �L$$��話������\$��� �Gl�$�Ѕ��L$ ���D$�����N ���ËL$d�    Y_^[��� �������U����j�hx�d�    P��SUVW�  3�P�D$0d�    ��~ ��   �N��Px�ҋN����@h�T$R�ЍL$�nQ���D$<    ������t'�L$�D$8���������ǋL$0d�    Y_^][��]Í�   R��b���؃���t�N��P|S�҅�u0S��b�����L$�D$8�����[���3��L$0d�    Y_^][��]�3�;��t$|?j ���r���������u	��;�~��#;�j���R���������Au�D$��;�~�D$S�qb�����L$�D$8����������D$�L$0d�    Y_^][��]������U����j�h��d�    P��hSVW�  3�P�D$xd�    ���|$ � �B  �O��Px�ҋ؃��-  ��   P�a���������t$�  �O��B|V�Ѕ���  �O��Rh�D$4P�ҍG ��P��Ǆ$�       �D$,���������   �D$4P����������   �U�K3���|D�N�B+�S���<�    �d$ �A�� �X؃� ���D��X��A��X��A��X�u܋t$�U;���+�+ʍ�����I ������X�u�V��`�����L$4Ǆ$�   �����e����   �L$xd�    Y_^[��]� j �L$8�p���j�ωD$(�s����T$$�����A��  j�L$8�G���j �ωD$(�J����D$$�������  3�V�ωt$(�+����}�T$��K��|7�J�Q�����uR�Q�����u;�����u7�Q����u2���C��� ;�~�;���k�������u��;�~��V����������;�C��I ����L$ j�\$0��虭���\$,����Au�L$�D$$�������;�D$$~t$ �\$$��j�΃��t$(�W����ߋT$R�_���D$$���x u�L$(Q���Q������p���3���|�I ���L$$���$�^�������;�~�T$ �z t)3��ۋ�|!���ǃ�����;��d��\�����\�~���3���������$    ���L$(���$辬������;�~������V��^�����L$4Ǆ$�   �����B���3��L$xd�    Y_^[��]� �����������V��~ tm�F�D$S�\$U�l$W�8SU���$������N���   ���$�ҋ���t.��t�E �����$������] ��t������$��������_][^� 3�^� ����j�h��d�    P��SV�  3�P�D$d�    ��3�9^��   �N��@h�T$R�ЍNQ�L$�\$(������t�N�D$,����   ���$�Ѕ����3���������;�t&��D$,���   �����$�Ћ���Bj�����ЍL$�D$$����������ËL$d�    Y^[��� �j�h�d�    P��SVW�  3�P�D$ d�    ���O��@h�T$R3��ЍOQ�L$�t$,�F�����t>�O�D$8�\$4��D$0���   ���$SP�ҋ������tS��tO� tI���FA �@����������t3�D$8�L$4��T$0���   ���$QR���Ћ���B���j�����ЍL$�D$(����������ƋL$ d�    Y_^[��� �����������̃y t�I�D$��T$���   ���$R��� 3�� �����̃y t�I�D$��T$���   ���$R��� 3�� ������j�hI�d�    P��SVW�  3�P�D$(d�    ��3ۉ\$3�9^t/�N��@h�T$R�ЍN�\$0Q�   �ȉ\$�Կ�����\$u�D$ ���D$0����t	�L$������|$ t �N����   �ЋL$(d�    Y_^[��$ËǋL$(d�    Y_^[��$������j�h��d�    P��SVW�  3�P�D$(d�    ��3ۉ\$3�9^t/�N��@h�T$R�ЍN�\$0Q�   �ȉ\$�������\$u�D$ ���D$0����t	�L$�1����|$ t �N����   �ЋL$(d�    Y_^[��$ËǋL$(d�    Y_^[��$������U������4SV��M$2���Wt�    �~ �,  �E�����$�����\$8�E�����$�u����\$0�EP�H5���E0�] �N���\$���E(�D$4�$P�D$DS�D$@P���\$�D$P    ��D$d���   �$W�҄��V  �D$(�����$�W����E�����E��z������A��   ������zi���������  ���D$0�D$$    ��4���D$8��4����������z��������{&������������   ��������A��   �����ًN�ۋ���E0���   ���\$�T$4�E(�$RS�T$@R���\$�$W�Є�tv�D$(�����$�w����E�E����������z��������{A������������   ��������z7���؋E$���M�t�T$$��_^[��]�0 ����������E�E������؋E;�t:�E0�M$�U���\$�E(�$QS��R���\$���$P��6��_^[��]�0 �����2���_^[��]�0 ����U����j�h��d�    P��hSVW�  3�P�D$xd�    ��~ ��
  �N��@h�T$$R��P�NǄ$�       蓻������L$$�؉�$�   ������t{�E��|s��
n��Rh�D$4P����j��Ǆ$�      ����� �]����Az��2ۍL$4��$�   �������t2��L$xd�    Y_^[��]�8 �EP�U2�����E�E8�U�N�9��(�\$ ���E0�\$�E(�\$�E �\$�E�$R�E���$�1����E�N���   ���$P�ҋL$xd�    Y_^[��]�8 �������V��W�~ ���r�����t�~ �����F��'���������_�   ^����������������D$SV��W�^ �����$�g���������;��������Au�D$$�ٙ��3�+�3Ƀ��������-��������������z�D$$�3�+�3҃��������|$$��t0�F��t�߄�uS�N迹����t���u������
��u�   �D$�����$�����~ ��   �T$(�N�\$����   U�l$ RW�|$,WUS���$�Ѕ��D$(��   �~ ��   �N��B4�Ѓ�|s�������3҃�|?�p������O��    �d$ �A��� �����Y��A����Y��A����Y��A����Y�u�;�}�d$ �׃�;����\��|����u��D$(]_^[� _��^3�[� ����j�h��d�    P�� SUVW�  3�P�D$4d�    ��u ��2��k�������   �}���Y�������   ��N�V�D$�F�L$�T$�D$ �L$DQ�L$�D$@    �����L$������tp�T$R�D$(P���2����L$$�D$<�������t?���%���L$$�T$(�D$,��L$0�W�T$�G�D$��T$ �O�L$�F�N�V��L$$�D$< �S����L$�D$<�����B����ËL$4d�    Y_^][��,� ���������U����j�h<�d�    P��(  SVW�  3�P��$8  d�    ��3�9F�;  �]S��$�   P�P����E�N��}���   ��$�   P���$WǄ$P      �҅��D$`��  �~ t����   ���ҋF �N$�V(�D$d�F,�L$h�T$l�D$p��Ƅ$@  t
S�L$h�s�����L$4j�L$h�r���j �L$h�D$@�c����T$<����\$��� �D$D�Pl�$�ҋG���8  ���/  ��Ph�L$<Q����j ��Ƅ$D  ����� �L$<�\$4Ƅ$@  �������Ph�L$tQ����j��Ƅ$D  �ܟ��� �L$t�\$<Ƅ$@  ������t:��躴���\$4����Au��訴���\$4�������\$<����z��������\$<�D$4����$�   �$P���5���D$<����$�   �$Q���5����$�   R���6����$�   P���w6��j������������!  ��$�   Q��$�   菨����u��$�   R��$�   �w�������   � u,��$�   Pj ���x����W��$�   Q��R���b����   �L$t�����L$<�ۥ����$�   P�L$x蚨��j ���q���ݔ$�   �D$t�L$t��Qj ���\$|݄$�   ��ݜ$�   ܌$�   ݜ$�   �t�����$�   R�L$@�C����G��P�������T$T�D$<�W�ɍL$<Q���\$@R�D$L�����\$L�L$T�\$T�"����L$dƄ$@   �������$�   Ǆ$@  ���������D$`��$8  d�    Y_^[��]� �������������̃y u3�ËI����   ������������j�hh�d�    P��SUVW�  3�P�D$$d�    ��3�3�9o��   �w��Ph�L$Q���ҍOP�l$0�l����L$���D$,�����������t6�GP�,0  ����t&��ȋBd�Ћ��t�U �GP���   ���Ѕ�t���L$<�D$4�Q�����$�w������   �����$�ҋ���t�\$<������$�������t�E �Pj���ҋƋL$$d�    Y_^][��� ����j�h��d�    P��SUVW�  3�P�D$$d�    ��3�3�9o��   �w��Ph�L$Q���ҍOP�l$0�\����L$���D$,�����������t6�GP�/  ����t&��ȋBd�Ћ��t�U �GP���   ���Ѕ�t���L$<�D$4�Q�����$�g������   �����$�ҋ���t�\$<������$�������t�E �Pj���ҋƋL$$d�    Y_^][��� ����j�h��d�    PQ�  3�P�D$d�    j0�83�����D$���D$    t���N����L$d�    Y���3��L$d�    Y���������������V�t$��th�����������t��^�3�^����������������j�h��d�    PQVW�  3�P�D$d�    ��j0�2�����D$���D$    t���������3����D$����tW���0����ƋL$d�    Y_^���������������VW�|$��t5h����������t%�t$��th����������tW�������_�^�_2�^�������������V�������D$t	V��3������^� ��j�h(�d�    P��SVW�  3�P�D$d�    ��|$(3�;��\$ t�^�b���N������N �����^�}��PS�҅�teS�D$0P�N 賜����tS�~S�L$0�b���� �����$������\$j�L$0�D���� �����$��������\$�L$<�D$ �$������3��Ή^����;��~t)�L$,�T$0���ĉ�L$D�P�T$H�H�ΉP�b�����D$,�L$0�T$4�F�D$8�N�V�F�V�F�N ��P�Q�P�@�Q�A�L$,�D$ �����f����L$d�    Y_^[��� �U����j�h��d�    P��   SVW�  3�P��$�   d�    ��t$$�~ ���D$(    �V������c  �^���D������Q  �Ej�����$�j������7  �E�����$�����T$,j�����$�?������  �E� 3�3���tP������������  �M���t#P������������  �U��M;��  �T$$�B�L$D�D$#�g����L$4Ǆ$�       �S����|$# Ƅ$�   ��t6j�[������\$�L$T�D$<�$�����D$,���$j ���1������4�D$,���$j �������L$T�$�ܨ��j���������\$�D$<�L$D�$輨���E�\$$���$�� j ���Ӗ�����L$t�$蔫��j��Ƅ$�   賖�����\$�L$d�E�$�m����L$DƄ$�   蜗�����b  �L$4苗�����Q  �L$d�z������@  �L$T�i������/  �L$$�Y����   ��Rh�D$tP����j �D$HP�L$|Ƅ$�   �L�����urƄ$�   �L$t������L$TƄ$�   �����L$dƄ$�   �����L$4Ƅ$�    �����L$DǄ$�   ��������3���$�   d�    Y_^[��]� j �L$8Q�L$|�Ƙ����Ƅ$�   �L$t�v����=�����u/j0�R-�����D$(��Ƅ$�   t	���h����3�Ƅ$�   ����u/j0�-�����D$(��Ƅ$�   t	���5����3�Ƅ$�   ���T$D�L$H���ĉ�T$\�H�L$`�P�HS��������T$4�L$8���ĉ�T$L�H�L$P�P�HS��������|$# t����   ���Ћ���   ���Ћj�L$h苔��j �L$h�D$,�|����L$(��Sl���\$��� �$�ҋj�L$X�V���j �L$X�D$,�G����L$(��Sl���\$��� �$�ҋE�8 u�0�E�8 u�8�D$(   �L$TƄ$�   ������L$dƄ$�   ������L$4Ƅ$�    �����L$DǄ$�   ���������D$(��$�   d�    Y_^[��]� ���������������j�h��d�    P��VW�  3�P�D$d�    ��|$,���F    t^��Ph�L$Q���ҋ���̉�P�Q�P�@�Q�AW���D$8    �Q����L$�D$$����������L$d�    Y_^��� �����N�_����N �W����F �L$d�    Y_^��� ���������������U����j�h �d�    P��hSVW�  3�P�D$xd�    �L$3��D$$%�\$(�\$,�\$0�};���$�   t9_|�_�u;�t9^|�^���L$ �y�����uD9\$0Ǆ$�   �����D$$%t�D$(;�tSP�L$,�%3��L$xd�    Y_^[��]� �D$9Xt��H��@h�T$4R�ЋL$ SQ�L$<Ƅ$�   �"�����u;�L$4��$�   �����L$$Ǆ$�   ������|��3��L$xd�    Y_^[��]� �L$ �T$4R�%������(  �D$�H����   VW�Ћ؃�}3�3�;�t9_t9G|�G;�t9F|�F3�;�t 9^t9F|�F;�t9G|�G3���   ;���   �L$8At;�t����6����t���7����tQ�L$����   �Ѕ�t?�G��~7��~�w�3����������V�P�N�H�V�P�N�H�V�u�P��tt�D$�x u�L$ �� P�Ŧ����tY3���~S�E�H��<�L$���$�`������;�|��-�L$���������t�E����   PW���ҋ؋�Pj���ҍL$4Ƅ$�    ������L$$Ǆ$�   �����#{���ËL$xd�    Y_^[��]� ������������V�t$��thx���������t��^�3�^���������������̸x������������VW����������~ t�N��P����~ t�N��P����~ t�N��P�����_^��������VW�|$��;���   W�
 ���N��t��Pj���F    �N��t��Pj���F    �N��t��Pj���F    �GP�|������t�O����P�g�����F�OQ�X������t�O�����P�C�����F�WR�-������t�O�ձ��P�-�����F_��^� ��j�h(�d�    PQVW�  3�P�D$d�    ��t$��w�N3�;ω|$t��Pj�҉~�N;�t��Pj�҉~�N;�t��Pj�҉~���D$��������L$d�    Y_^����V��~ t>�~ t8�N��Pj �҅�t(�N��P4�҃�thdyhHyjeh(y�L�����3�^� �N��Pj �҅�t�~ tM�N��Pj �҅�tԋN��P4�vW�ҋ���P4����;�_th�xhHyjnh(y������3�^� �   ^� ������̋D$h�yP��#����� �����������V���Pj �҅�tS�FW�|$P����������t;3�9N��Q����!������t$�N��tQ���c�������t�VR���Q�����_^� ��������̃�SV��N3�;�Wt	��Pj�ҋN;�t	��Pj�ҋN;ˉ^�^t	��Pj�ҋ|$�D$P�ω^�\$�Y�����t)�D$;�t!P������;ÉFu�L$;�t	��Bj�ЍL$Q�ω\$�\$������;�tA9\$t;�T$R�������;�t+�L$;�t#Q�m����;ÉFu�L$;�t	��Pj��3�;É\$tH�D$P��������;�t4�D$;�t,P�*����;ÉFu�L$;�t	��Bj��_^3�[��� ��_^[��� ������̃y t
�I��P4��3��������������̃y t
�I��@8��3�� �����������VW�|$W�������������~ t�N��PDW��_^� _3�^� �������������̃y t
�I��@P��3�� �����������j�hi�d�    P��VW�  3�P�D$ d�    ���D$    �t$0���D$(    �~���� �D$(    �D$   t.�O��@h�T$R�Ћ��P�V�H�N�P�L$�V�����ƋL$ d�    Y_^�� � ���̃y t
�I��Px��3��������������̃y t
�I��@|��3�� ����������̃y t�I����   ��3�����������̃y t$�T$�D$�I����   R�T$R���$��� 3�� �V��~ tD�FP�������t4�NQ�������t$�N�D$����   ���$�Ѕ�t	�   ^� 3�^� �������������V��~ t5�FP�^������t%�D$�D$�N����   ���$P�D$P��^� 3�^� �����������̋AP����������� �����������V��~ t�~ t�N����   �҅�u��^���^������̃y t�y t�I����   ��3������V��~ Wt4�N����   �ҋ���t�~ t�N����   �ҋ��������_^Ë�3�������_^�����h�yh�yh�  h(y�{����3�� ���������������j�h��d�    PQVW�  3�P�D$d�    j���������t$3�;��|$t*���|
����w�~�~�~�ƋL$d�    Y_^���3��L$d�    Y_^��������j�h��d�    PQSVW�  3�P�D$d�    ��j�C�������t$3�;��|$t����	����w�~�~�~�3�;��D$����tS�������ƋL$d�    Y_^[����������������VW�|$��t5hx���������t%�t$��thx���������tW���V���_�^�_2�^�������������V�������D$t	V�{ ������^� ��U�������  SVW����$�   �   �I ��艍������y�$�  �   ��I ���i�������y�L$X�X�����P4���҉D$���������3�;��  �E ;��L$,�L$0�L$4t#� �Ё��  ���T$,����%�   �T$4�D$09Ots9Otn�G�U�0�L$,QR��$�   ���   �Ռ���E�]�OP�jS���$�Ѕ��D$��  ��3���~Hܔ$�   ��ܜ$�   ��A��z��Az�   �'��_^[��]� �   ���Az�   �	�   ��؋O�1�T$0RP��$�  �ư   �C���݄$�   �OP�jS���\$݄$�   �$�Ѕ��D$��  �E ��t$�L$0�T$4�����   ʋT$,������  ʉ�|$݄$�  ���u�~
݄$�  �^��~
݄$�  �^�E�������D$�q  ݄$�   ��$  P�\$$݄$�   ����$�   �T$$�$Q�����D$0��P��$�   R��$�  P����$�   �$Q������������� ���T$X�@�T$`�@�T$h���~�^��؃�~�^���t$����  ݄$   ��$P  �\$@R݄$  ���\$D��$�   �D$$���T$|�D$,���\$\�$P�[����D$0����P��$�   �L$Q��$@  R����$�   �$P�*����D$h��P��$�  Q��$0  R����$�  �$P������D$X��P��$\  Q��$   R����$�  �$P�Ԍ���D$h��P��$|  Q��$  R����$�  �$P詌�������ϋ�����ȋ�����������躋��� �T$X�@�T$`�@���T$h���~�^��؃�~�^���t$���{  ݄$  ��$�  �\$xQ݄$$  ��ݜ$�   ��$�  �D$,����\$T�D$|�L$$�$R�����D$X�D$(��P�ɍ�$d  P��$�  ��Q����$�  �$R�Ћ���D$`�L$8��P��$T  �L$$P��$�  Q����$�  �$R蝋���D$p�L$@��P��$�  P��$�  Q����$�   �$R�n����D$@�����P��$�   �L$TP��$p  Q����$�   �$R�9����D$p�L$H���D$XP��$d  P��$`  Q�L$L����$�  ������$R�����݄$�   �L$x��P��$  P��$P  Q����$�  �$R�Ȋ��݄$�   ��P��$  P��$@  Q����$�  �$R蚊��݄$�   ��P��$�  P��$0  Q����$�  �$R�l�������蒉����苉����脉�����}������v������o������h������a���� ���T$X�@�T$`�@���~�^��؃�~�^��؋D$���|(���D$    ������~�V��~�V���u��؋D$_^[��]� ����̸h������������j�h�d�    PQSVW�  3�P�D$d�    ��t$�q���~���D$    �<z� ���   ���D$�w���H+���\$�����D$,�$hhY� ����� ݞ�   ǆ�      �ƋL$d�    Y_^[�������j�hC�d�    PQSUVW�  3�P�D$d�    �ى\$�����{���D$     �<z�� ���   ���D$ ��~���D$,�t$(�&   ��] �D$4ݛ�   ǃ�      �ËL$d�    Y_^][��� ��������j�hs�d�    PQSUVW�  3�P�D$d�    �ى\$�l$(U�;���{���D$     �<z�C ���   �D$ �#~���u�&   󥋅�   ���   ���   ���   ���   ���   ���   ���   ���   ���   �ËL$d�    Y_^][��� �����j�h��d�    PQV�  3�P�D$d�    ��t$�<z���   �D$   �_����N�D$ � ���D$�����s ���L$d�    Y^������k ���   ������V��L$�FPh�   Q��m  ���   RjP�m  �ư   VjP�m  ��$^� �����SU�l$��;�tSVWU����u�{�&   󥋅�   ���   ���   ���   ���   ���   ���   ���   ���   _���   ^]��[� ����������U������4SVW���w���( �؅��  �D$P��� �D$�} ��   �U�����z�����D$�R����z�Z����D$(�M�����Au�����D$0�Q����Au�Y��؃��   ��   �D$ �R����z�Z����D$8�Q����Au^�Y�L$������_^[��]� �E�M��D$�X�D$(��D$0�Y���   ~$�D$ �X�D$8�Y�L$�^�����_^[��]� �؍L$�H���_^��[��]� �������������VW�|$W�������������W�N� _��^� ����������VW�����   ���?|����u;�|$��t,j���{�����$j ���{�����$h@{W�����_3�^� �O�x ��u�D$��th{P�a����_3�^� _�   ^� ������������̃�0SVW�����   j���z�����$j ���z���t$H���$h�{V��������{��h�{V�������_S������݇�   ���$h�{V��������� ���$h�tV������D$P�������L$$Q���5��h�tV������T$R���[��h�tV�p�����D$$P���A��h�&V�V���������_^[��0� ���VW�|$j ��j���-������t8�FP���B������t&���   Q���3������t���   R���1����_^� ��������̃�VW�|$��D$P�L$Q���D$    �D$    ��������tc�|$uZ�VR���;2������t&���   P�����������t���   Q�����������   ��t��t_ǆ�      ^��� 3�_^��� ���D$V�D$3���W������z*�����\$���   �$�R����Ͼ   �&���_��^� �ً�������_��^� �������������VW�|$�G�����w)9��   S�t�����3Ƀ��������   ��[_^� _2�^� Q�D$���   ����   �P���   ���   �P�$    �HY� �������������VW���   j ���w���|$j����w���_���x��_��^� �������������̋D$��S��t�D$����$P���   ����   W�|$��tV�s�&   �^��_t��Bj ����[� ���   u�D$�D$���$P��6��� W�|$��tV�q�    �^�   _� ���D$�D$���$P���i' ��� ��̃�� �������V��N� ��t���   �fz�����_����   ^���������U����j�h��d�    P��h  SVW�  3�P��$x  d�    ��$�   �}��3ۍ��   S���Pv���\$\j���Cv���\$\����A��  �D$l�^P���5
 ��Ǆ$�      ��v���\$\����v���|$\�L$lǄ$�  �����\$|������L$\�\$lQ����	 �D$L�E�����$Ǆ$�     �v���L$L���$�u���L$\�\$LǄ$�  �����T����D$L�b �\$T�D$L�>c �D$T������4������AtL������4������{=����������{������zL�������������������z�0'�-���)�������������������������z�0'�����܎�   �F8P���\$`��$   �~ ܎�   �T$h�$R�~���D$d��P��$�   PW����$�   �$Q�`~����P��$�   R���}}�����v}��݄$�   �}�݄$�   �_���   u
݄$�   �_�E����   �]�D$l��ۉD$L�L$|�F8P���\$x��$�   �D$`�D$h���\$`�T$h�$P��}���D$d��P��$   Q�F P����$@  �$R�}��������|��� ݔ$�   ��@ݔ$�   �@ݔ$�   �D$l����������_���   u���_��؃l$L�Q����ظ   ��$x  d�    Y_^[��]� �Ë�$x  d�    Y_^[��]� ��������U����j�h!�d�    P��   SVW�  3�P��$�   d�    �ى\$P�}���D$H    �t�������D$L�<  ����   �����$�2s���\$T�G�����$�s���\$\�D$d��P���� �D$T���L$l�$Ǆ$�       �r���\$T�D$\���L$l�$�r�����D$T������;����AuR�����\$��$�   �$�'�������̉�P�Q�P�@�Q�A��Ƅ$�   �D$X   �u ��t������2��D$HǄ$�       t	�L$t������t���W�V�G�F�O�N�t$L�3��L$P�����L$dǄ$�   �����}����Ƌ�$�   d�    Y_^[��]� ���U����j�h��d�    P��   SVW�  3�P��$�   d�    �����   �҅�t2���$�   d�    Y_^[��]� �D$,P�L$HQ��2��A����}j ���%q���\$D����zj ���q���\$D�j���q���\$,����Auj����p���\$,���t���������Rh�D$TP���ҋ؍D$4�~P��Ǆ$�       �� �D$(�D$D�����$Ƅ$�   ��p���L$(���$�p���L$4�\$LƄ$�    �2����L$TǄ$�   ����������Rh�D$dP���ҋ؍D$TP��Ǆ$�      �G �D$(�D$,�����$Ƅ$�   �jp���L$(���$�p���L$T�\$4Ƅ$�   趾���L$dǄ$�   ����袾���D$L�H+�T$4������   �L$T�\$4Q���� �؋�Rh�D$dP��Ǆ$�      �҉D$(�D$4�����$Ƅ$�   ��o���L$(���$�o���L$d�\$,Ƅ$�   �����L$TǄ$�   �����	�������D$4���\$��$�   �D$\�$���������̉�P�Q�P�@�Q�A��Ǆ$�      �� �L$tǄ$�   ����覽���D$,��Bl���\$���D$T�$�а��$�   d�    Y_^[��]� ̋�Pj �����������������������j�h��d�    P��   SVW�  3�P��$�   d�    ��$�   �D$P�L$Q���D$    �D$    ����������   �|$��   �L$�� �T$R��Ǆ$�       �t������D$P�N�T  ��t&���   Q�����������t���   R�����������   ��t��t
ǆ�      �L$Ǆ$�   ����� �ǋ�$�   d�    Y_^[�Ĝ   � ���������������j�h��d�    PQ�  3�P�D$d�    h�   �%�����D$���D$    t���;����L$d�    Y���3��L$d�    Y������������V�t$��thh���������t��^�3�^����������������j�h�d�    PQVW�  3�P�D$d�    ��h�   ������D$���D$    t���������3����D$����tW���M����ƋL$d�    Y_^������������VW�|$��t5hh����
�����t%�t$��thh����������tW�������_�^�_2�^�������������V�������D$t	V��������^� ��U������4SV��W�~��2�� ����   �E�Ơ   �����$��k���H+���\$(� �D$(P�����$�U j���lk��� �Ej ���\$,�Zk���D$(��� �L$@�\$�E�$�������P�V�H�N�P�L$0�V�������_^[��]� _^��[��]� �����U����j�ha�d�    P��h  SVW�  3�P��$x  d�    �ٍ{��� ��t3���$x  d�    Y_^[��]� 3����   t���]����D�  �L$d�q���L$L�q����Ph�L$4Q����j�ȉ�$�  �Yj��� �L$4�\$,Ǆ$�  ���������D$,VV�D$TP�L$pQ�����$�R����L$L�x����$�   ��  �UR�D$PP�L$lQ��$�   Ǆ$�     ��  ��;ƉD$,t��$�   �  �&   ��$�   ��  ��Rh�D$4P����j��Ƅ$�  �i��� ����$�   �$P��������L$4Ƅ$�  �G����MQ��$�   �'����\$4���|	 ��;�\$4����A��   ���pp��P�T$8R��$�   �^r����K �P�s �V�H�N�P�V�H�N�P�ΉV�w��V���)	 P��$�   P�y����S8�P�K8�Q�P�Q�P�Q�P�Q�@���A�Mw���H+�����$�� �D$,   ��$�   Ǆ$�  ������  �t$,���@����Ƌ�$x  d�    Y_^[��]� ������U����j�h��d�    P��h  SVW�  3�P��$x  d�    �ٍ{��� ��t3���$x  d�    Y_^[��]� 3����   t���]����D��  �L$L�o���L$|�o����Ph�L$4Q����V�ȉ�$�  �g��� �L$4�\$,Ǆ$�  �����p����D$,VV��$�   P�L$XQ�����$������$�   �t�  �UR��$�   P�L$TQ��$�   Ǆ$�     ���  ��;ƉD$,t�&   ��$�   ��  ��Rh�D$4P����V��Ƅ$�  �g��� ���D$l�$P���<����L$4Ƅ$�  軵���L$dQ�M螅���\$4���� ��;�\$4����A��   ����m��P�T$8R�L$l��o����K �P�s �V�H�N�P�V�H�N�P�ΉV�u��V��� P��$�   P�%w����S8�P�K8�Q�P�Q�P�Q�P�Q�@���A��t���H+�����$�d  �D$,   ��$�   Ǆ$�  �����5�  �t$,�������Ƌ�$x  d�    Y_^[��]� U����j�h&�d�    P��   SVW�  3�P��$�   d�    ���|$L��Ph�L$TQ���ҍD$d3�P�O��$�   ��  �ES���L$`�$Ƅ$�   ��g�����L$du;Ƅ$�    �$����L$TǄ$�   ��������3���$�   d�    Y_^[��]� Q�L$X�{���E��u���L$\�$�fe�����L$l�$�e��S���L$p�$�Gg����u	�L$d�y����U�3���t�M;t�P�����������t֋��r����U���tP�����؃���t����S�����u?h�   �u������D$P��Ƅ$�   tW�������Ƅ$�   ���3�Ƅ$�   ���;�tW���4�����u?h�   �&������D$P��Ƅ$�   tW������Ƅ$�   ���3�Ƅ$�   ���;�tW�������;��L$T��   j ��c���E���\$��$�   � �$�x���P���   ��Ƅ$�   �ЍL$t��Ƅ$�   �o�������   j�L$X�c��� ���\$��$�   �E�$�Qx���Ƅ$�   ���   j�Yc��� ���\$��$�   �E�$�x���P���   ��Ƅ$�   �ЍL$t��Ƅ$�   ������thj �L$X�c���E���\$��$�   � �$��w���Ƅ$�   ��P���   �ЍL$t��Ƅ$�   蔱����t�E�8 u�0�E�8 u>��:�M�9 u9t$Lt��t��Bj���ЋM�9 u9\$Lt��t��Bj���ЍL$dƄ$�    �/����L$TǄ$�   ���������ǋ�$�   d�    Y_^[��]� �U����j�h[�d�    P��l  VW�  3�P��$x  d�    ����  ��u3���$x  d�    Y_^��]Ë��i��� ݜ$�   ���@ݜ$�   �@ݜ$�   ��  �D$|�\$,P�����  j ��$�   Ǆ$�      �a��� j�\$@��$�   �ua��� ��$�   �\$lQ�����  ���I�  ��t	��$�   ���$  R�����  ��L$T�P�T$X�H�L$\�P�T$`�H�L$d�P�T$h��$4  �D$8   ��I ���)h���� �l$8y��8�D$,��������Az	�ظ   �� 8����A�   {�   �< ���O�L$8�C  ����$�   ��$4  R�w  �j���D$,�Xe����$$  ���D$D�$P�7 P��$X  �Zj���D$,�8'����$�  �T$L�D$D�$Q��� P��$x  �&j���D$,��|����$  ���D$D�$R�� P��$�  ��i���D$,��$����$4  ���D$D�$P� P��$�  ��i���D$,��|����$�  �D$D�$Q���s P��$�  �i���D$,�@'����$�  ���D$D�$R�C P��$�  �fi���D$,��|����$\  �D$D�$P��� P��$  �6i���L$TQ��$8  �%i���D$D�\$,�	  �i���D$,�8'����$  ���D$D�$P�� P��$X  ��h���D$,��$����$t  �T$L�D$D�$Q��� P��$x  �h���D$,�@'����$�  ���D$D�$R�\ P��$�  �h���D$TP��$�  �nh���D$D�\$,�U��$�   Q��$8  �Ph���D$,��$����$�  ���D$D�$R�� P��$X  � h���D$TP��$x  �h���D$,��$�J ����   ;����D$<ݔ$�   ݜ$�   ~u݄$�   ��$\  ��݄$�   ��݄$�   ���D$,��������@���@;��X����@��X��@����X����P����P�̴݄   ��ݔ��   ݜ��   |������؃��ًL$8���D$lݔ��   ݜ��   �|  ����$T  �����    ���F�L$t�T$,Q�����T$P��T$H�T$X��{�$�a} ���������D{���X<����Az�D$t�`�����D$L�T$<����D{�L$,�����D$D��$�   �NR���T$H�T$X��{�$��| ���������D{���X<����Az݄$�   �`�����D$L�T$<����D{	�L$,�^����F��$�   �L$DP���T$H�T$X��{�$�| ���������D{���X<����Az݄$�   �`�����D$L�T$<����D{	�L$,�^��؃�@��������L$8��؋u3҃���3��K�C   �C   �������S���C ��P���n����D$8��P���ϓ��3�9t$8~L��$<  V���(���G��}���Xu�G�X��G�X�G�X݄��   �K����� ;t$8|��S�D$l�D$8�L$|��Ǆ$�  �����٩���   ��$x  d�    Y_^��]����������������S�\$j�����������[� ������U����j�h��d�    P���   SVW�  3�P��$�   d�    ��$�   � ���3ۋΉ�$   ��  ���  �};���   �D$TP���q�  S�L$XƄ$  �?Z���E� S�L$X���\$P�*Z��� �L$T����|�\$L����uKS�Z��� �L$T���$   �Ǩ����$�   Ǆ$   ������������$�   d�    Y_^[��]� j�Y���E� j�L$X���\$P�Y��� �L$T����|�\$L����uj�y����ES���$��[����uA�L$T��$   �6�����$�   Ǆ$   �����O���2���$�   d�    Y_^[��]� ��$�   Q���F�����t��L$d�I`���E����$�   �$R��$�   �<�����L$d�P�T$h�H�L$l�P�T$p�H�L$t�P�ΉT$x��_��P�L$h�ba���D$dP��$�   ��`���L$|Q����_�����N3��P�8i���\$T���T$dR��$�   �`���D$|P���_�����-3��P�i���D$T���W �\$DS�L$X�MX���D$D� ���5H+�$��F ����S�L$X��$�l$H�\$H�X��� �\$D����Atj�L$X�X��� �\$D����z?j�L$X��W��S�L$X����W��� ��L$T��$�]����AuS�j�W��� �\$D�L$T�|X����|����Au{�D$D���L$\�$��W���\$L�E���L$\�$��W���p&�����H���Au�T$L����z�ڍL$T�����6�����������z�\$L����Auj�L$X�������D$D���������������U����j�h��d�    P��(  SVW�  3�P��$8  d�    ���w�  ����  �}����  �D$DP�����  j�L$HǄ$D      �V��� ��j �L$H�\$8�V��� ��j �D$8�L$H�h,�\$@�rV���E� �D$<������uJ��N����u?j �L$H�HV��� ��L$DǄ$@  ����� ������$8  d�    Y_^[��]� ��j�L$H�	V��� �E���D$<������uP��N��������AzAj�؍L$H��U��� �L$D�Ǆ$@  ����菤�����$8  d�    Y_^[��]� ��j ���L$P�$��W����t:��$�   ����j��$�   ��Ƅ$D  �:���������u;Ƅ$@   �T����L$DǄ$@  ��������2���$8  d�    Y_^[��]� �q���j �L$H�D$\�U��� ��$�   �\$t�0\�����)\��P�L$`Qj ��$�   ��x������$�   �$R��$�   ��������]��P��$�   ��\����$�   P�L$`�\���L$\Q����[�����C/��P�-e���\$D����$�   R�L$`�\���D$\P���[�����"/��P��d���D$D����R �\$43�3�9\$X�  ���g[��P��$�   Q�SR��$�   �.x�����D$l�$P��$�   �G������0]��P��$�   �\����$�   Q�L$`��[���T$\R���[�����.��P�id���\$D����$�   P�L$`��[���L$\Q����Z�����^.��P�8d���D$D���6R �D$4������z���
���H+���D$t�T$t���\$4�]����AtS��$�   ���yw���;|$X�������$�   �{��v��;�|+j�L$H�S��� �U��$�   �Ƅ$@   ��������W��$�   �w�����$S��$�   ��v������$�   �$�g����$�   Ƅ$@  �	L  ��$�   PS��$�   Ƅ$H  �\�����u4��$�   Ƅ$@  ��Y  ��$�   Ƅ$@  �@�����$�   ������$  �������$�  �l+������Ƅ$@  �kY��PW��$  �=�����$�  Ƅ$@  ������$  Q��$�   �d  �E3���R �\$4��$    V��$�   ��R  � �L$4V��$�   �\$@�R  �D$<�����`�\�T|��D$d�����D$l���D$\�������T$4���������T$<����;����A�Z  ������������Az�   �3�hd}h<}h�  h }P�F���D$H���P& �D$\�d$d�����D$<�����T$4��������At��������z-����������$��������������������Au���T$4�
����������h<������Az�}����Az	�   ���3�h�|h<}h�  h }P��E��������D$4������������z~���ك���$�   �$�P���U��$�   �Ƅ$@  ��W  ��$�   Ƅ$@  ������$�   Ƅ$@   �)����������������������������D{!�������w�����������A�u������p������������c������������������j�h+�d�    P��   SUVW�  3�P��$�   d�    ��$�   3�;��\$trV�L$�����W�L$��$�   �5�����t!݄$�   ��$�   S���$P�L$(�����؍L$Ǆ$�   �����l����Ë�$�   d�    Y_^][���   � ���   ���1P����tэn����  ��tË��   ��$�   Q����������t3�+j�Ͼ   ��N�����$j ����N���Ul�����$�ҋ��v����D$�m����������U����j�h`�d�    P��hSVW�  3�P�D$xd�    ���D$$�wP����  ���E�Ǡ   �����$Ǆ$�       �N�������$�SN���\$�L$$Ǆ$�   ���������D$�L$Q�����$�E����T$4R������  �D$�����$Ǆ$�      �:N�������$��M���E�L$4�Ǆ$�   ����脜���ËL$xd�    Y_^[��]� �������������U����j�h��d�    P��hSVW�  3�P�D$xd�    ���D$$�wP���s�  �D$�E���   �����$Ǆ$�       �M���L$���$�?M���L$$�\$Ǆ$�   �����כ���D$�L$Q�����$���������tP�T$4R�����  �D$�����$Ǆ$�      �"M�������$��L���E�L$4�Ǆ$�   �����l�����E�M��ǋL$xd�    Y_^[��]� �����������j�h��d�    PQV�  3�P�D$d�    h�   �4��������t$3�;��D$t���J�����{�ƋL$d�    Y^����V�t$��th@����۰����t��^�3�^���������������̸@������������V���H�����}��^��������������̋D$VP���3�����}��^� ������̋D$VP���3�����^� ���������������}鵵�������U����j�h��d�    P��SVW�  3�P�D$ d�    ��t$�L$������P4���D$(    �ҋ؃��U�M����T�P�L$���������Q��j V�<��# ���} t]�E� �U��@�^�@�E�^��� ��@�_�@�_�} t,������{�A�Z����{�A�Z����z�E    �E�L$��R8PWV�҃��D$~(��E��F�X�F�X�E���G�X�G�X�"������M�Q�E�P�Q�X��؍L$�D$(����������D$�L$ d�    Y_^[��]� �������������U������   S�ً�P4VW3��҃����ww�E��wo�}��wg;�u�F_^[��]� ����L$H�$�m���3�V�L$D�Q�����9uu���;�u�M���������|Ӌ�RD�D$@P����_^[��]� _��^[��]� ���������������   ܜ$�   V������Dz��ܜ$�   ����Dz�   ^�Ā   � �L$����݄$�   ��$�   ����ĉ�Q�P�Q�P�Q�P�Q�I�P�H��$�   ����ĉ�Q�P�Q�P�Q�P�Q�I�P�H���\$�L$D݄$�   �$�"�����RD�D$P����^�Ā   � ������������V�D$����������Dz�ظ   ^� �D$�L$PQ��4 ���$�D$��5 �����$�����^� �́�   VW��$�   �����W����t_�   ^�Ā   � �L$�[���W�L$������PD�L$Q����_^�Ā   � �������̋D$P�&����   � ��������������V�t$��� ��^� �������������̋���D$�����P����H����P����H����P2�� ��V����}�b����D$t	V���������^� ������������j�h)�d�    PQVW�  3�P�D$d�    ���D$    �t$ ���D$    �����j �FPV���D$$    �D$   �2�����u���g����ƋL$d�    Y_^��� ̋D$P�D$�PRP������ ����������j�h`�d�    P��@SUVW�  3�P�D$Td�    ��t$h���|$dt���Y����u	3��������\$l����   ������$���������   j�L$������L$$�D$\    �����j �D$@P�L$,Q���D$h�P�����t#�T$R�L$(����SVW�L$ ��C  ��t�   �L$$�D$\ �K����|$  �D$\�����D$�$t-�D$��t%j P�L$��$�V�GPW���������t�   �����L$Td�    Y_^][��L� ������������V�t$��th0����۩����t��^�3�^���������������̸0������������j�h��d�    PQV�  3�P�D$d�    ��t$��~�N�D$    �������D$�����Ӯ���L$d�    Y^�����V��N�E�����~ �~  |f�~4 vf���    u	�   ^� 3�^� ����������́�   �  3ĉ�$�   V��$�   Wj��j����������   �G P�����������   �OQ���p�������   h�   �T$j R�� 3�����@�O4}f�f�TD������@|�D$Pj@���������t>�OQ���j�����t/�WR���Z�����t�G�����$�������t��$W���'�����$�   _^3����� �Ą   � ����������̸   � �������̃�`�  3ĉD$\SW�|$l2ۅ���   f�? ��   Uj �`!���t^Vj\�D$j P�
 �t$8��3ɋ�+��f��tf������� |�j j h@u�L$QU�D$;� ��^u�Uj �\!]_��[�L$\3�� ��`ËL$d_��[3��� ��`�����SUV��F3�;�}3�;��   t���   ��  8^��:��   t���   ��  8^��:��   t���   ��  ���   W2ҋſ    ���    ��`���f9tf������u�:�_tU�������������   ��  ^][���VW�|$��t5h0����z�����t%�t$��th0����b�����tW���ֳ��_�^�_2�^�������������V�������D$t	V�;�������^� ��SV��W�N�s����؅�u��7�F �|$PhTW����Sh@W�����N4Qh(W�����VRhW�����FPh�~W�{����NQh�~W�k�����@�F�$h�~W�W�����_^[� ��������������SW��h�   �_4j S� �D$����tRV�H3��G6���    �Q�f��t7f�P��Q�f��t*f��f��tf�P�Qf��tf�P��������@|�^j@���   j P�O ����Ǉ      ����f�; _��[� ��������������̋D$;At��}3��Aǁ      �o���� ������������V��W�N�������~3��^�F�  �F �F �F �����F$�F(�F,h�   P�F0�F4P� j\���   j Wǆ      � ��hh���   Ɔ�   ����_^���������������̊D$8At�����Aǁ      ����� �������������j�h��d�    PQV�  3�P�D$d�    ��t$�S����N�D$    ��~�������D$������ƋL$d�    Y^�����������������U������$  �  3ĉ�$   SV�uW���|$�t$����3��D$�D$�D$P�L$Q�_ ����������������   �|$��   S�������؄���   ��W��������؄���   ��$�   Rj@���"����؄���   �    ��$�   �|$ �t$�D$ P���D$@   fǄ$�     �����|$��   �|$�L$Q���y����؄�ts�T$R�������D$P���[����؄�tU�|$ ��Q���5����VR��������؄�t4�|$|-��$V���B������h�h�h�   ht�0����2ۋ�$,  _^��[3�� ��]� ������j�h��d�    PQ�  3�P�D$d�    h  ��������D$���D$    t�������L$d�    Y���3��L$d�    Y������������j�h�d�    PQVW�  3�P�D$d�    ��h  �Q������D$���D$    t���G������3����D$����tW��荮���ƋL$d�    Y_^�����������̸ ������������VW�|$W����l�����   ���   ���   ���   ���   ���   ���   ���   �R���   ���   ���   P�ҋ��   ���   ���   ���   ݇�   ݞ�   ݇�   ݞ�   ݇�   ݞ�   ݇�   ݞ�   ��   ��   ��  ��  ��  ��  ݇  ݞ  ��  ��  ��  ���  �P��   �H��$  �P_��(  ��^� �������m����x��������SV�t$Wjj��h � @���'q���؄���   ���   P�������؄���   ���   Q�������؄�to���   R���c����؄�t[���   P���O����؄�tG݇�   �����$������؄�t.݇�   �����$�����؄�t݇�   �����$�����؋��;�����}��td݇  ܏�   �
��tR݇�   �����$�m����؄�t9��   Q��������؄�t$��  R�������؄�t��  P���@����؋��Ǘ����}��tE���
��t=݇  �����$�����؄�t$��  Q���O����؄�t��  W���+����؋��"�����u	_^��[� _^��[� �����������̃�SV�t$3�W�D$�D$���D$P�L$Qh � @���T���|$��t2��   ����   ���   R���޾���؄���   ���   P�������؄�tt���   Q��蒼���؄�t`���   R���~����؄�tL���   P��������؄�t8���   Q�������؄�t$���   R���Ҽ���؄�t���   P��込���؃|$|<��t8��   Q���s����؄�t$��  R��������؄�t��  P��苼���؃|$|(��t$��  Q���`����؄�t��  R��輻���؃|$|��t��  W��������؋�������u_^��[��� _^��[��� �����������̋D$h�P�q������   � ������V�t$��th����;�����t��^�3�^���������������̸������������j�h}�d�    PQV�  3�P�D$d�    ��t$�$����   �D$   ��������   �D$��������   �D$�������   �D$�����N�D$ �������D$���������L$d�    Y^�����SV��3��F�����F�F�FhP��N3ۉF�h�����$�V �   �V(h�7�荎�   �V0�FP�ɉ^T�^8�^X�8'�^\�^@�^`�Fh�Fd�VH�Fl�����^p�^x�H'���   ݞ�   ���   ���   ���   �����h�7���   �����h`����   �����h\����   ������ݞ�   ���   �艞�   ���   ݞ�   ���   ^[�V��N�e�����~�~ |	�   ^� 3�^� ������������VW���O��������u��7�G�|$Ph��W�����Vhh�W�������_^� �̃�VW�������|$�D$P�L$Q���D$    �D$    �����|$����  ���&  �VR��许�������  �FP��舽��������   �N Q������������   �V(R�������������   �F0P������������   �N8Q���и��������   �V@R��躸��������   �FPP����������tz�NTQ����������th�VXR����������tV�F\P���޷������tD�N`Q���̷������t2�VhR��躷������t �FdP��訷������t�NlQ��薷�����|$|��t�VHR���������|$�'  ���  �FpP������������   ���   Q���3���������   ���   R������������   �FxP���t���������   ���   Q��苷��������   ���   R����������tz���   P���Ͷ������te���   Q��踶������tP���   R��裶������t;���   P���~�������t&���   Q���i�������t���   R���d������|$|��t�FP���k������|$|��t���   Q��迶�����|$|^��tZ���   R��裶������tE���   P�����������t0���   Q���I�������t���   V���4���_��^��� 3�_^��� ��������������̋D$�Al� ������VW�|$��t5h ���芖����t%�t$��th ����r�����tW������_�^�_2�^�������������Q��SV��ݖ�   h�   ݞ�   3���h�   ݖ�   h�   �L$ݞ�   ���   ǆ�      ��   ��  �ٰ����D$ݞ  ��  3�9��   ��  ~��$    ���   ���;��   |�^[Y���������VW�|$��t5h���蚕����t%�t$��th���肕����tW��薣��_�^�_2�^�������������j�h��d�    PQV�  3�P�D$d�    ��t$�Ӓ���N�D$    �$��������   �D$��������   �D$��������   �D$��������   �D$��������D$�a����ƋL$d�    Y^�����������������V�������D$t	V��������^� ��j�h&�d�    P��SUVW�  3�P�D$(d�    ��t$�n_��3퍾�   ����l$0��H�o�o�o�   ��  �\$0�����D$P� ��z�����N�P�V�H�N�P�V� 0�F�0�N�0�V �0�^(�F$�G�B   ;�}@9_~�_��G�RSP����;ŉGt�O;�}��+�R�UQ�� ���_��o�o9_|�_�`/���   �d/���   �h/���   �l/���   �`/��  �d/��   �h/��$  �l/��(  ��������ƋL$(d�    Y_^][�� �j�hX�d�    PQSVW�  3�P�D$d�    ���|$���3�9��   ���   �\$��Ht�F;�tSP����H�^�^�^���D$������^���L$d�    Y_^[�������������j�h��d�    PQ�  3�P�D$d�    h�   �e������D$���D$    t��������L$d�    Y���3��L$d�    Y������������j�h��d�    PQVW�  3�P�D$d�    ��h�   ��������D$���D$    t���g������3����D$����tW���͟���ƋL$d�    Y_^�����������̃�V�D$��P� ��ێ��P���c�������th ����a�����t݆  ^�����^��������������j�h��d�    PQ�  3�P�D$d�    h0  �%������D$���D$    t���k����L$d�    Y���3��L$d�    Y������������j�h�d�    PQVW�  3�P�D$d�    ��h0  �������D$���D$    t����������3����D$����tW�������ƋL$d�    Y_^������������V���8����D$t	V�K�������^� �̃�W����t:V�D$P� ��v���P�����������th ����������t��Bj����^���u���_���U������8��V�u�\$4W����������}���'����\$8jj���h��������R  �GP��蒿�������<  �OQ���,��������&  �G ���L$@���$����������  �G(���L$@���$�����������  �G0���L$@���$����������  �G8���L$@���$����������  �G@���L$@���$����������  �WPR���˾�������u  �GTP��赾�������_  �OXQ��蟾�������I  �W\R��艾�������3  �G`P���s��������  �OhQ���]��������  �WdR���G���������  �GlP���1���������  �GH���L$@���$貿��������  �Gp�����$藿��������  ���   Q������������  ���   R���u��������o  �GxP������������X  ݇�   �����$�0��������:  ���   Q���w��������!  ���   R���^��������  ���   P���E���������   ���   Q���,���������   ���   R�������������   ���   P������������   ���   Q������������   �WR��軾������ty݇�   ���L$@���$�M�������t[݇�   ���L$@���$�/�������t=���   P���z�������t(���   Q����������t���   R��������_^��]� ���V�t$��th ����+�����t��^�3�^���������������̸ ������������V�t$��th���������t��^�3�^���������������̸������������V�t$��thЖ��請����t��^�3�^���������������̸Ж�����������VW�|$W���B����G�F�O�N�W�V�G�F�O�W�NR�N������� W�N �����_��^� �����V�t$��th����������t��^�3�^���������������̸�������������j�hS�d�    PQV�  3�P�D$d�    ��t$�c����N�D$    �T�蝹���N �D$萹��3��F�F�F�F�F�����ƋL$d�    Y^�����������j�h��d�    PQV�  3�P�D$d�    ��t$�T��N �D$   �B����N�D$ �5������D$����膏���L$d�    Y^��������V���P4W�ҋ|$Ph�W襻����P8������Ph؁W荻����P<������Ph��W�u�����PD������Ph��W�]�����_^� �����V������3��F$�F(�F,����^����SV��F$��Wt�N,��t��u	P��������F$    �N(��t�F,��t��u	Q�������F(    �~���F,    �"����^ ������3��F�F�F�F���F�����̷��_^��[�·����V��~$ t'�~( t!��P4�҅�~��P8���҅�~	���^� �D$S2ۅ�thT�P�Z�������[^� ���������������j�h��d�    PQV�  3�P�D$d�    ��t$���D$    ��������D$����������L$d�    Y^�������̋A$��t�@�3���̋A$��t�@�3���̋Q$3���t �V�r�P4���ƃ���������^������̋A$��t�@�3��̋A$��t�@�3����SUV���P@W�ҋ؋F$��t2�H �|�(��t'��t#�l$��|��P8����;�}�����_^][� _^]3�[� ��������������̃�43�SUV�L$3��D$�D$�D$ �D$$�D$(�D$,�D$0�D$4�D$8�D$<�����l$D�D$P�͉t$�t$������؄��%  �L$�T$�L$R���ߥ���؄��  �D$�L$Q�͉D$ ������؄���  �T$�D$P�͉T$$�����؄���  f�L$�T$f�L$$R�������؄���  f�D$�L$Q��f�D$*�c����؄���  �T$�D$P�͉T$,�E����؄��m  �t$�L$Q�͉t$0�'����؄��O  �T$�D$P�͉T$4�	����؄��1  �L$�T$�L$4R�������؄��  W�|$�D$P�͉|$@�̤���؄���   �L$�T�,R�L$D�D$ (   �����������tj,j W��� ���(   ���D$�x$u_^2�]��[��4� �
   �t$�@,   �3�9t$<~a��t]�|$�G$�L�(Q��肢���؄�t;�W$�D�)P���m����؄�t&�O$�T�*R���X����؄�t�G$�L�+Q���C����؃�;t$<|��T$0��v!��t�L$�A$�t$<�D�(P�A(R���1�����_^]��[��4� ��̃�4SUV3��ىt$�=����l$D3��D$�D$�D$ �D$$�D$(�D$,�D$0�D$4�D$8�D$<�D$P�͉t$�t$�k������W  �L$�T$�L$R���O������;  �D$�L$Q�͉D$ �3������  �T$�D$P�͉T$$�w������  f�L$�T$f�L$$R���Y�������  f�D$�L$Q��f�D$*�ۢ������  �T$�D$P�͉T$,迢������  �t$�L$Q�͉t$0裢������  �T$�D$P�͉T$4臢�����s  �L$�T$�L$4R���k������W  W�|$�D$P�͉|$@�N������9  �L$�T�,R�L$D�D$ (   �\���������tj,j W�i� ���(   ���{$��   �C,   �
   �t$�|$0���C$� (   v�K$�T$<�D�(�C(�L$HQ���D$L    ��  ����   �t$<�D$H��;�t�>;�thP�h,�h  �t�S$�L$Q��(RP���<�  ��tk��vg9t$Hua�D$HP���D$L    �J�  ��tI�D$H;�u#�S$�L$Q�L$@�T�(RP�����  _^][��4� h�h,�h  ĥ������2�_^][��4� ���SUV��F$3�;�Wt�~,uP�U������n$�~�ωn(�n,�n0�ܯ���^ ���ү��3��F�F�F�F���F����膰��_^]��[�{�������������̃y$ u�D$��th�P�7�����3�� �   � �������V�t$Wj ��j����������tF�G P����������t4�O0Q���)�������t"j����������t�W$�G(RP�����  ��_^� ����������̃�VW���D$    ������|$�D$P�L$Q���D$    �D$    藶��������   �|$��   �V R���D$�����~�������t�F0P���|����L$Q���p�������tQ�L$�� StO��uA�^(S���?�  ����t/���vP�l������F$�F,   �F$��T$RPQ�����  ��[_^��� �^(S����������t���vP�"������F$�F,   �V$�RP���7���[_��^��� _3�^��� �j�h��d�    PQVW�  3�P�D$d�    j0覲�������t$3�;��|$t*���������~$�~(�~,�ƋL$d�    Y_^���3��L$d�    Y_^��������j�h�d�    PQVW�  3�P�D$d�    j4�&��������t$3�;��|$t-����������~$�~(�~,�~0�ƋL$d�    Y_^���3��L$d�    Y_^�����VW�|$W��肉���G�F�O�N�W�V�G�F�O�W�NR�N�8����G P�N �,����O$�N$�W(�V(�G,�F,�O0_�N0��^� �������������VW�|$��t5hЖ���:~����t%�t$��thЖ���"~����tW���V���_�^�_2�^�������������j�h;�d�    PQVW�  3�P�D$d�    j0���������t$3�;��|$t*��������~$�~(�~,�|��ƋL$d�    Y_^���3��L$d�    Y_^��������V�������D$t	V�{�������^� ��V��������D$t	V�[�������^� ��QSU�l$��;���   ����U�������E$����   �@ V�4�    �E �PDW�͉t$�҉D$�D0,P����������tj,j W�,� ���(   ���{$t_�D$���C,   �u$�
   �~�M$�S$P��(Q��(R��� ���T$��~F�C$��t�H �3ɍD�(�C(�m(��RtUP��� ��_^]��[Y� j P�� ��_^]��[Y� _^]�C(    ��[Y� �������������VW�|$����au����W��u�����_��^� �G���_��^� ���������������V���|��b����D$t	V��������^� ������������j�hh�d�    P��SVW�  3�P�D$d�    �ً|$(�D$P�L$Q���D$    �D$    �S�������tv�|$uo�L$(�L����T$(R���D$$    �8�������u�L$(�H����W���n������D$(P�K �ΰ���L$(�D$ ���������ƋL$d�    Y_^[��� 3��L$d�    Y_^[��� ��������������̃�,�ыB$2Ʌ��$t�R(��t�x v�H �L�(;�����SUVW��t.���@ �
   �|$�L$��,�    �BD�Ћ����D$u.�*3�3�3��D$�D$�D$ �D$$�D$(�D$,�D$0�D$4�D$8��t$@P���6������   �L$Q���"������  �T$R����������   �D$ P���Z�������   �L$"Q���F�������   �T$$R���ҩ������   �D$(P��辩������   �L$,Q��誩������   �T$0R��薩������   �D$4P��肩����tp�L$8Q���r�����t`��t9�T$�B$���/t��(PQ��� �  _^][��,� 3�PQ����  _^][��,� �\$�C$��(PU�����  ��t�K(QW�����  _^][��,� ����j�h��d�    PQV�  3�P�D$d�    ��t$����D$    ��������D$�����F����L$d�    Y^��������j�h��d�    PQSVW�  3�P�D$d�    ��j0胫�������t$3�;��|$t���i������~$�~(�~,�3�;��D$����tS��������ƋL$d�    Y_^[����������������VW�|$��t5h�����w����t%�t$��th�����w����tW������_�^�_2�^�������������j�h��d�    PQSVW�  3�P�D$d�    ��j4裪�������t$3�;��|$t����������~$�~(�~,�~0�3�;��D$����tS�������ƋL$d�    Y_^[�������������VW�|$��t5h�����w����t%�t$��th�����w����tW������_�^�_2�^������������̋D$P������� VW�|$j ��j���}�������t�F P���[�������tW���������_^� ����V�������D$t	V苫������^� ��j�h+�d�    PQSVW�  3�P�D$d�    ��j0�S��������t$3�;��|$t���9����~$�~(�~,�|��3�;��D$����tS��������ƋL$d�    Y_^[���������������̋L$W�|$���j  ���b  ���D$V�  U�����I �����4Ux3Ҋ��������f3���3������4Ux3Ҋ��A�������f3���3������4Ux3Ҋ��A�����f3���3������4Ux3Ҋ��A�f3���3������4Ux3Ҋ��A�f3���3������4Ux3Ҋ��A�f3���3������4Ux3Ҋ��A�f3���3������4Ux3Ҋ��A�f3���3ƃ��������]��t0���    �����4Ux3Ҋ�f�����f3���3ƅ�u�^_�f�D$_���������������W�|$���)  �D$���  ��V�t$����   U������3ց��   ������3�x�3с��   ��3�x�P3с��   ����3�x�P3у����   ��3�x�P3у����   ��3�x�P3у����   ��3�x�P��3с��   ��3�x�P��3с��   ��3�x���������*���]��t$��I �3΁��   ��34�x������u��֋�^_ËD$_����̋A�L$��� ���V��W3��~�~�~9~|�~�F ;�tP�L������~ �F,;ǉ~$�~(�~,t��    �pP�'�����;���u�_^������������SU�iV2�;iWu�Y��Y�Q(�t$�|$+�+���t6��|2�Q;�}+��|';�}#;�t3҅�~������������;Q|�_^][� ����������U������4�Q;QSVW�L$ u�A��A��I3��\$8;щD$�t$$�T$,~�L$,3�9t$,�D$�c  �L$�]�L$��d$ �D$�L$��	�1�H��D$��+����L$(��   �|$���G��0��������Au�ىL$��؋G��0��������Au�A�ىD$��؋�0��������Au�A�ىD$��؋G�0��������Au�A�ىD$��؃��B���;��{���;�}&�D$���0��������Au�ىL$��؃�;�|��D$8�L$������At��u�T$8�]����A�J  �D$$9L$td�|$ ;Wu�G��G�$�D$0�D$+�+ϋ|$0��t(��|$;�} ��|;�};�t���T$0�����D$0���D$�ËL$�����T$����40ƋT$ ��PP���T$@���X��B+����$P�h   ��L$D�L$4�|$<����Q;�}p�T$���0����T$0��������]����Au@���I+L$�D2PP�D$ ��D2P�����$Q�.   ��L$H�L$8��������؋Q��;�|��D$(�D$��;D$,�D$�������؋E��t�D$8��D$$_^[��]� ����S�YW�y;�~_2�[� V�t$;���   ;���   ��;�U�l$ }�D$�D� ��������At��;�|���;yu�A�D$�]��^_2�[� �I�L$�D$$���;�t�D� �؍s���|3+ލ<�+萋D$���WR�T�RS�Z  �,/�����������}�]^_�[� ^_2�[� ����V��~ ���t%�F��tj P����F    �F    �F    ^�����������V��~ ���t%�F��tj P����F    �F    �F    �D$t	V��������^� ������SV��F 3�;���tP�W������^ �F,;É^$�^(�^,tW�xP�7�����;���u�_��9^���t�F;�tSP������^�^�^^[���QSUW��2������|$���  �|$ ��   9}V�u}W���[����} ��   ;~�~�L$���3Ҹ   ���;�&��}�u�   �u�|$�";�}k����;�|�ߋu�u�|$��|$;�}�ߋ��|$��   R�����H�H�8�U,�P�E,�@��C�����t�L$����у��V����u�D$+Ã����D$��D$�L$^_�E�M]�[Y� ^_]��[Y� _]��[Y� �������V���X����D$t	V�[�������^� ��j�h[�d�    PQV�  3�P�D$d�    ��t$3����F�F�F�F���F�F�F�L$�D$�F �F$�F(�F,�D$ PQ���F����ƋL$d�    Y^��� ̋D$�T$P�D$R�QP�AR�QP�A�	RPQ�I]���� � ��̋�3ɉ�H�H�H�H�H����������̋D$V��3Ʌ���3�W�|$��#�9T$���3������V��#ǅɉF~��3����F����N�NPQ觸������ɉF_2�^� �V��t��u�S�^��|�~�;�|�v��~��;�}[_2�^� [��_��^� �����U�����M��t��SVW�  ����$輛������   �L$8�����L$P�����]�D$4    �|$4 �Et
� 3��\$8��@3��\$8��E��t�@3��\$@��@ 3��\$@��E��t�@��@(�L$8�\$HQ�M�T$lR������L$P�P�T$T�H�L$X�P�T$\�H�L$`�Pj �D$TP�ˉT$l��T����t1����|������o����D$4�����D$4�<����_^[��]�2�_^[��]ËMj Q�M��X��_^[��]������������̃�0SU�l$@��VW�|$D��t�������u3�\$L����   ������$�c�����umV�D$P���2���U�L$Q����Y����V�T$,R��������L$�P�T$�H�L$�P�T$�H�L$ �Pj�D$P�ωT$,�Y��_^]�[��0� UV���Y��j��V���Y��_^]�[��0� U����j�h��d�    P���   SVW�  3�P��$�   d�    ��}��tv������$膙����uc�H+���$V�L$8�̢  �E�MWPQ�L$8Ǆ$      ��
  �L$,��Ǆ$   �����i�  �Ë�$�   d�    Y_^[��]� �]�ۋ}t�������u3��FX���\$�FP�$���܎�   �\$4�FH�\$�FX�$����܎�   �\$,�FP�\$�FH�$����܎�   ������D$$����   �������Au��������W����Au�_����F�D$���G������Au���_����F�W ����Au�_ ����F���W����z�_����F�W(����Au2�_(�/�����_�F�D$�����_�F�_ �F���_�F�_(��ذ��$�   d�    Y_^[��]� ��������̃��(�����������U����j�h��d�    P���   SVW�  3�P��$�   d�    ��}���]t�������u	3����NP���~ �(  ��$�   �O���}��Ǆ$       ��  ������$�3������s  �L$L�R���FP�L$hQ���������$�   �P��$�   �x��$�   �X��$�   �X��$�   �@��$�   ��$�   ��$�   �   9~��$�   ��$�   ��$�   ��$�   ��$�   �0  �   �I �F�P�L$hQ�M�]���� �T$L�@�T$T�@�T$\݄$�   ������Au��ݜ$�   �݄$�   ������z��ݜ$�   ���݄$�   ������Au	ݜ$�   �݄$�   ������z	ݜ$�   ���݄$�   ������Au	ݜ$�   �݄$�   ������z	ݜ$�   ��؃���;~�*����P�T$dR���LP��� ݜ$�   �L$d�@ݜ$�   �@ݜ$�   �@ݜ$�   �@ ݜ$�   �@(ݜ$�   �8N���M��$�   P�xQ����$�   �   Ǆ$   �����N��3�������$�   d�    Y_^[��]� ������������̋A��t�I�L$��� 3�� �����̃y t�A��t�Q�T$��� ��� ��������������SV��F����I  �L$���=  ;N�4  �V��W�<ЋD$������  �$����L$���PQW�� ���~ th����׊�_^[� �~ �T$t���   QRW�r� ��_^��[� ��U�.��������D{�4�3Ʌ�]~��+�����Ƀ��X�;|���_^��[� �~ �T$t.���3Ʌ�~��+�����Ƀ��X�;|���_^��[� ����QRW��� ��_^��[� �~ �6t���L$��    PQW�� ��_^��[� _2�^��[� ^2�[� �I ��#���׺������������SV��FW�|$3�;�~H�N;�u"��    P�*�����;ÉFu'�^_^��[� ;�~��    RQ�c�����;ÉFtى~_^�[� �������������̋�3ɉ�H�H�H�H�H�H�H�����V��NW�|$;�}:�F��t��t/��    QP����������    R膮�����F���#ǉF�~ _��^� ������������D$���$��������tt�D$��$����D{a��������Dz�ذËL$���T$�D$V�t$����+ʃ�t)W�<�    �ҋ�t� ���Ƀ����X�u���Ƀ�u�_�ذ��^���2�����U�����E��4SVW���$�f���������  �E(���$�M���������  �E������������D��  �E(��������D��  �U����  �M$;M��  ;�u��������D��  ��������z��������A�o  ��������Au��������Au��2���_^[��]���;�~�ɉU$�]�M�ыM$�](����؋}�]�u�������Ӄ����T$@���\$8�$�d���������  �D$0���$�J���������  �����D$8��������D��  ���D$0��������D��  ��������z��������A��  ��������Au��������Au��2���_^[��]��ڋE���M$tB;�t>�}(+ȉL$(���u���D$(������� �T$(�E�t$8�\$8�E��� �|$8�\$0�.;��E�����T$0t�E(�����E$������ ��������\$(�D$(���$�K���������   ���\$(������   �D$0���$� ���������   �D$0��$����D��   ��M��������D{?��+���~'�хۋ�t����ʃ����^�u��    ���u�����ǃ��؍4����D$(��������D{VWQS���$����������E���}$�M������E(��_^[��]�������_^2�[��]���������V��FW3�;�t9~~	P�Ȫ�����~�~�~�>�~�~_^��j�h��d�    P��  SUVW�  3�P��$�  d�    ����  3ۄ�t9��$�  ;�t����$������t��$�  ��$�  SPQ���"����  9�$�  t��$�  �h����u��$�  ��$�  �F����$�   �   ��I ��������� ��y�L$0�9���L$0�T$\��$�   Q�͉�$�  �T$P�D$\蒜������   ��$�  ;�t������$�P�����u
V�L$4�<���\$,�D$@�T$D�\$8�l$<�L$P�|$X�p����;�Ƅ$�  �\$�l$�D$ �L$$�|$(}i��    �D$�D$L�D�������Au6��$�  ��$�  �D$$j Q�L$(RWPQUS�OM���� ��tǄ$�     �T$D|$�����;�|$(|�3�9�$�  �\$X�\$L�L$0��Ǆ$�  �����of���Ë�$�  d�    Y_^][���  � ̃�������������̃��x�����������j�h(�d�    P��0SUVW�  3�P�D$Dd�    ���t$X���l$Tt���	����u	3�����D��� ��   �D$P���������\$\�D$L    t(S�L$QU���������t�L$�D$L�����mD����[��t)������$膋����uSVU�O������t�   ��T$R���G�����������L$�D$L�����D��3������L$Dd�    Y_^][��<� ��������U����j�hX�d�    P��   SVW�  3�P��$�   d�    ��t$ �]3�9}t���g����u�}�D$TP���ԭ����$�   �}����  ������$裊������  W�L$XQS��������t.�L$TǄ$�   �����DC�����$�   d�    Y_^[��]� �F���D$�>  �VR�L$(�n����D$$P�L$@Q��������L$T�P�T$X�p�t$\�x�|$`�X�\$d�@�D$h��$�   �D$���L$l�T$p�t$t�|$x�\$|��   �]�   �x���T$ �B�P�L$(������L$$Q�T$@R��茈��� �T$$�@�T$,�@�T$4�D$T������Au���\$T��D$l������z���\$l����D$\������Au�\$\��D$t������z�\$t����D$d������Au�\$d��D$|������z�\$|��؃����@����]�} u8�D$T����D$\�[�D$d�[�D$l�[�D$t�[ �D$|�[(�g�����E��L$TQ����D���} �L$T��Ǆ$�   �����xA���Ë�$�   d�    Y_^[��]� �������������̃� W��� �|$�D  U�o��V�7�t$�+  �G;��   ���  ;�Su	�^�\$��D$�؋���P���������l$ ��   ��F���������������҉D$,�t$$�T$�G��t�O�͍<��3��L$����|$,�|$�|K�q���T���+��ݍD�����B�� �X(�� ���D �X �B(�X�B �Xu܋l$ �|$�t$$�T$��|�׍�+���������}�T$�D$�|$(�Ã���l$ �t$$�N����\$�؉_�G   [� ^]��_�� �V��FW3�;�t9~~	P�X������~�~�~�~�>�~�~�~_^������������QW��� �  �O��V�7��  �G����  ����  �WS�_;�U��   ;��^����P��������O�G�W���Íi���D����   ��O���L$x�O��t�W�_���\$Ӎ��3����3ۃ��L��|2�V�������    ��� �X �� ���A�X�A�X�A�Xu�;�}��+�����X����u��l$y����l����؋G����]�G   � [�w�G^��_Y�;֋��^����P��������O�W�G���Ӄ���D���L$��   ��o��x}�O��t�W�_���\$Ӎ��3����3ۃ��L��|2�V�������    ��� �X �� ���A�X�A�X�A�Xu�;�}��+�����X����u���y��l$�p����؋G����]�w�G�G   [� ^��_Y������SVW�|$����|{�F;�}t�\$��|l;�}h�D$��$����D{U���$�D�������tE�D$ ��$����D{2���$�!�������t"���D$�����D$ ��z������Au������_^2�[� ��������Au��������Au_��^��2�[� ��;�u��������Dz�;�~�\$�ǋ��\$ �������W��������\$����DzS������\$ ����Dz_^�[� ���2����D$ �F�N�V���$S�D$ ���$WP�QRP�������(_^[� ���������������V��~ W�|$u)���W`����Dz�Wh����Dz�_p����D{	��������F�N�VWP�FQ�RPQ�0  ��_^� ��������j�h��d�    P��(SUVW�  3�P�D$<d�    ��~u'�F�8 t�ȋD$T�	��R<P�D$TP�D$TP���  �l$P��t�L$L�9 ����u3�L$L�z;���F����   �P�L$�6��3�9~�D$D    ~H�d$ �N�<� ��t0��T$$R����P�L$�~����N���D$$P�~���P�L$�d�����;~|��\$T�T$LSUR�L$ �X�����t�   3�9~~-�F�<� t�ȋ���D$L�R<SUP�҄�t�   ��;~|Ӄ|$  �D$D�����D$�$t�D$��tj P�L$��$3������L$<d�    Y_^][��4� �̃��x����������̋D$��u�D$� �L$�	Ã�u�D$�L$�@�I� �	��Ã�u�D$�L$�@�I� �	���@�I��Ã�u%�D$�L$�@�I� �	���@�I���@�I��Å���t�L$�T$����	��������u���̋D$��~"�D$�L$�T$����Ƀ������Y�u���������V�t$��~,�D$�D$�L$�T$����Ƀ��������A��X�u���^���������̋D$��~"�D$�L$�T$����Ƀ������Y�u����������D$���D$���D$����������4����������t>������������A{5��������Au�������������4��������t�   �����������3��L$��t������������������U������tSV�uWV��������\$�}W��������\$W�������j ���\$�D$4�\$�D$,�$�!����؃��ۉ\$u�M�����M ������_^[��]�W�D$$VP��������L$ �s����T$�������\$��4����z�M������M ����3�_^[��]ËM�A�E�O�]�G�U �I���F�H���F�H�����I��O���F�����H���[�G�	��I�M����H���F����[�G�H�G�H���F�I���F�I�����H� �O���F�	����I���Z�G���H����I���F�	�L$ QS���Z�����t$���T$D�$R������D$(��P�D$TP���L$x�$Q���>�����������u ��H�K�P�S�H�K�P�L$ �S�@QV�C�����t$���T$t�$R�s����D$(��P�D$TP���L$H�$Q���������������\$��H�N�P�V�H�N�P�V�@_�F^��[��]����������������D$�D$������z��2��ȅ���   �D$������z�����������Au����������������������4����S��4��������u
����$��ًD$������t���������ًD$ ��t�������؋���������U������   SV�uW��������\$ �}W��������\$(�������j ���\$�D$D�\$�D$<�$� �������tW�D$LVP��������y  �L$0�L����L$`�C����L$H�:����E��t$��t����u�\$ �0'��0'�T$ ��0'�\$ ��M�T$(Q����$�   �$R�����D$0�]��P��$�   PS����$�   �$Q�`������������ �T$0S�@���T$D��$�   �@�T$L���N���N���\$T���N������\$\����N���\$d�D$4�$R������D$0�M��P��$�   PQ����$�   �$R��������������� �T$0�@�T$8�@�T$@�G���G�����\$`��G�D$`��P�L$|Q��L$P�\$p�G������\$x������M ��P�Q�P�Q�P�Q�P�Q�@�A����_^��[��]���������U������xV�uW��3������T$0��������Dzx�u�؋�������������zG���D$@�$P���q�����M��P�Q�P�Q�P�Q�P�Q�@�A�M������_^��]ËM�������M������_^��]Ã��L$@�$Q��������u�}��H�N�P�V�H�N�P�V�@V�L$<Q�ωF������������D$0��V�����T$D�\$<�$R�5�����P�D$TP���U����D$0P���L$t�$Q������M��P�Q�P�Q�P�Q�P���Q�@_�A�   ^��]�������������̋L$�V�D$�t$�у�������z�����^�������u������A�F��   ��^��Q����z3���^��T������u�F���^��AW�3�����Dz�D���������D{��D��������Dz�D����������D{�G;�}Z�>��������z#�D����������Dz4�D����������D{��!�D���������Dz�D���������D{�W;�|�����_^����̃�V�t$��W��   �|$����   ����   ����   ���>�L$��   ����   ��u��+_^��Ã�u��'_^��Ë�%  �yH���@t%�O�QV�~����\$W���V�p����D$��_^��Ë�����~%�W�RV�P����\$W���V�B����D$��_^���;�~+΋���H�����_^��������D$_^�����_^�����_^������������V�t$��W|>�|$��|5�T$��|,�|$$ t%�|$ t���L$;�|�D$ ;�|;���;�}_3�^���;�|�_�   ^����Q�D$��SUV~%�T$�ҍHu�ȋl$ ;�|�t$��|�\$$��u^]2�[YÅ�t����~|W�<�    W�>�������������D$�D$    ~G�,���D$WSP�D� WUS�<� �L$0WQU�0� �L$H�T$4��    �+��$�+�;։T$|��T$R������_^]�[Y����������Q3�9D$$�$u/�D$ �L$�T$jP�D$Q�L$ R�T$P�D$QRP������� Y�V3�9D$~XS�\$$U�l$$W�|$0�D$$���͍ϋL$R�T$SPQR��������t��u�D$   ��;t$ |ƋD$_][^Y�_]3�[^Y��QSV�t$���	  �\$����   �D$����   �T$����   �L$ ����   ;���   ;���   ;���   ����   U3��|{W��{�������,�    �d$ ���\$�����D$������\$�����D$������\$�����D$������\$�����D$��ƃ�u��t$_;�}%��+ݍd$ ���\$�����D$��ƃ�u�]^�[Y�^�[Y�^2�[Y���SV�t$����   �\$����   �D$����   �T$����   �L$����   ;���   ;���   ;���   ����   U3��|\W���{�������,�    �I �����������������������������������ƃ�uËt$_;�}���+݋���������ƃ�u�]^�[�^�[�^2�[�������������̋L$��3�����   �D$����   �T$S�U�l$�Vҋ�L$0�T$�T$,W�t$,�D$3ۃ���|_�t$(���}��������    ���    �����������������������������������ƃ�u�;�}"�|$(�����+���������ǃ�u�t$,t$�l$�t$,�[���_^][�   �����������̋D$��SUVW�~%�|$���Hu�ȋl$ ;�|�t$��|�L$$��u_^]2�[ËT$(��t��u_^]�[Å��I  �����  ����   �<�    ����J �A�J(���A�J0�����J8���A�JH��J@���A�JP�����JX����J`�A�Jh���A�Jp�����Jx���A�J��
���A�J�����J������Y�Y��υ��s���_^]��[Í�    ��I ����J �A�J(���A�J8����J`�A�Jh���A�Jx���A�J��
���A�J������Y�Yȅ�u�_^]��[Í�    �����J`�A�Jx����
�A�J����Yȅ�u�_^]��[Ã�����<�    �  ����   ����J`�A�Jh���A�Jp���Bx��������Dz��2��������J �A�J(���A�J0���B8�A�JH��J@���A�JP���BX�A�J��
���A�J���B��������Y���Yυ��o���_��^��]��[�����J`�A�Jh���Bx��������Dz��2��������J �A�J(���B8�A�J��
���B������Yυ�u�_��^��]��[�����J`�Bx��������Dz��2��������
�B���υ�u�_��^��]��[������������̋D$��SUVW�~%�|$���Hu�ȋl$ ;�|�t$��|�L$$��u_^]2�[ËT$(��t��u_^]�[Å��I  �����  ����   �<�    �B(���I�B �	���B0�I�����J8���BH�I�B@�	���BP�I�����JX���B`�	�A�Jh���Bp�I���Bx�����A�J��
���A�J�����J������Y�Y��υ��s���_^]��[Í�    ��I �B(���I�B �	���B8�I���B`�	�A�Jh���Bx�I���A�J��
���B�I������Y�Yȅ�u�_^]��[Í�    ��Bx���I�B`�	����
�A�J����Yȅ�u�_^]��[Ã�����<�    �  ����   �B`���	�A�Jh���Bp�I���Bx��������Dz��2�������B(�I�B �	���B0�I���B8�BH�I�B@�	���BP�I���BX�A�J��
���A�J���B��������Y���Yυ��o���_��^��]��[��B`���	�A�Jh���Bx��������Dz��2�������B(�I�B �	���B8�A�J��
���B������Yυ�u�_��^��]��[��B`���	�Bx��������Dz��2��������
�B���υ�u�_��^��]��[�������������QV�t$$3�W3�9D$�D$~b�D$ S�\$0��    U�l$,�L$0���T$$�D$�L$SVURPQ��������u
�D$    ���u�D$   t$0��;|$ |��D$][_^Y������V�t$��W~�|$;�|�T$��|�D$��u_3�^ËL$��t����   ����   ���4�    t[�d$ � ���I �@�I(���@�I0��� �I@�@�IH���@�IP��� �	�@�I���@�I������X�Xƅ�u�_�B^�� ���I �@�I(��� �	�@�I����Xƅ�u�_�B^Í4�    ��I � ���	�ƅ�u�_�   ^����������V�t$����   �T$��L$�D$����   ����   ����   ������������Dz��������Dzq3�������������D��   ��;�X<������؋ƃ�����   �������B���������������A{���������������������t���������2�^�����;�X<������؋ƃ���tD������������������A{���������������������t���2���^��۰��^������ٰ��^���������������SV�t$����   �\$��|{�L$��U�l$�Eu��W�|$ ;�|Y������Ǎ�RVQU�z�������t>�|$~��u_]^�[Ð�|$ �D$�<�WVPU���I�������t�ۋ�u�_]^�[�_]^2�[�^2�[���������̋T$��ҋL$VW�|$t������D{	�����4�������ҋt$t��������D{�4����3҅�~w�X<��;����̃��F���������������������z��������������At?��������{H����4����������At#��������At��;�|�������_3���^���������_�ڃ����^�����_�ڸ   ��^���U������t��S�]V�uW3��}�|$(uq��l9}~g�؃����$�&�������tN������������D{@�E �������$���������t$�M ������������D{���D$'�T$0��������D$' ���T$0���T$8���;����9}�ʉ|$,�\$@���\$H�T$h�T$p�T$x�T$P�T$X�\$`�3  ���+  �M �U�EQSRP������������   �|$' ��   �D$0�$���\$@����A��   �D$8�M �$���\$H����A��   �|$( u�|$(V�T$lSR聬 �D$t�4�} V�D$`WPݜ$�   ݄$�   �4ݜ$�   ݄$�   �4ݜ$�   �B� �D$h�4>�E�L$hQ��$�   Rj P�\$x݄$�   �4>ݜ$�   ݄$�   �4>ݜ$�   �-�����(�����#|$(�M�E �U�ˍЋD$,��;E�M �D$,�������_^[��]��W�|$3���~XV�t$��~N�L$$��tF9D$(t�D$����t$ �����D$ ����|$��RPQ�L$P�D$ VPQ�����������^_�����������������D$��������DzS�����D$��������Dz(�D$ �؋L$���\$����D�������  �������ًT$ �|$�D$�����������D$��������DzV�����D$��������Dz�L$ �؋T$����   ������������z�D$�L$ �3��ËT$�ɋD$ ��3�����D$��������DzA���������T$���/� �L$ ����T$����Au�T$����   ËD$�����3���������H'��������������4������u�������������A��   ��V� 5�t$ �������������Dz�L$$����   ^�����菢 ��$�D$�L$$�������������D$�������D$��������z	������t������Au"������Az���������������   �^�������������������������t������������������tŸ   ^��ܸ   ���������^���������ϡ �D$����������$��������z�����D$���D$������������Dz�T$ �ًD$���������   ���������Au����� 5���T$��������   ������A��   ��������������������������������t]������������������������tP��������z	������{:��������AuA������Au<�ًL$ ���D$�T$��   ����������������������������������؋D$�ɋL$ �3������U������E4�M0��U,��E8��M����t��S�AV��W��3�3�����Au�ٍ_����A��������Au	�ٻ   ��؋u���������Au�ٿ   3�����F��������Au�   �ً�����F��������Au�   �ٍ_��؋U���������Au�ٿ   3�����B��������Au�   �ٍ_�����B��������Au�   �ً������������Dz��3���_^[��]Ã����T$�\$��   ��tU��E�E�D$ �A�D$$�A�D$(�A�D$,�A�I�D$0��L$4�N�D$@�F�L$D�N�D$H�F�L$L�N��   ��E$�D$ �E�B�T$X�D$$�E�B�D$(�B�D$,�B�R�D$0��T$4�V�D$@�F�T$D�V�D$H�F�T$L�V�D$P��T$T�Q�D$`�A�T$d�Q�D$h�A�I�T$l�   ��E�D$ �E�F�D$$�F�D$(�F�D$,�F�D$0�F�D$4��D$@�A�D$D�A�D$H�A�D$L�A�I�L$T�T$X�J�E$�D$P��L$d�J�D$`�B�L$l�J�D$h�B���\$x�D$p�L$ttM���}0�  �D$ �E,�D$0�U4�\$ �U,���\$0�D$@�D$P�\$@�T$P�D$`�D$p�\$`�\$p�D$H�D�D$ �E,�D$(�M0�]4�\$ �M,�\$(���D$@�D$H�\$@�T$H�D$`�D$h�\$`�\$h�D$P�����t$ �D$(���T$(�D$0���T$0�������T$8�D$@����������D{q���������T$H���������T$P�����������\$X�����D$`����������D{<�����D$h�\$h�����D$p�T$p�����D$x�\$x� �D$P�]4�D$H�Z�������������D$p����3���3�����������Au�ٍN����D$h��������Au�پ   3��������������Au�   �ً��������������Dz�ٸ   ������������_^[��]������D$������z�\$��D$������Au�\$��؅�t2�̋��\$(�]0�ʋ��\$0�E4���\$H�\$P�D$h���\$h���\$p�
���������م�t
�L$h�T$H��L$H�T$h����q����������I�Y�D$(����������D{����Ƀ��D$0�\$0�I�D$8�\$8����������������D{����Ƀ��������I�B�Z��������������Dz�ظ   ��_^[��]������D$������z�\$��D$������Au�\$����:����A�����������D{�
������D$0����������D{�
�D$8����D$8���U,�t�D$x��D$X�
�D$X��D$x��E8�D$_�t$^[��   ��]�������̋L$�A�T$��R�T$�ЋAR�Ѓ���������������̃� S�\$4���e  W�|$0���W  U�l$@���I  ��u]�    _[�� �3҅ۋË�t�����Յ�u�L$D3��|$0�D$ �D$$�D$�D$(�D$8V�D$$�L$(��u�T$ Rh �jSW�������   ����L$�����t�l�����(�L$�T$����l��(�T$��T�tt�t	;�L$wZs�L����Q�R�T$0�����D$$}�����T$�QR�T$0����}���L$�t$���t6��s;�D$$v��L$�T$�,����^����\$@�/�l$D�ۋ�t��$    �3��������ɉF�u�^]_[�� �����̋L$��W�|$(����������Dz	��2�_��ËT$ ��U��l$(�BV���Ņ�t����Ƀ����^�u�����`  �ɍ�    �4:����S�T$����t��+��(���Ƀ����@��X�u�l$0�|$,�  �����2�ȋ���t!����Ƀ����N��������@��X�u߃|$,������   ��+��D$ ����    +����   �9l$,�|$4��   �D$0�AȍωD$�L$�3ۅ�L$~s�l$��I �T$SR�u����D$ �+D$$�L$0�������D$��t������������F��^�u�l$�؍�    +��D$ ������;�|��|$4�T$T$��;l$,�l���[^]�_�����[^]�_������������������U������DSV�uW�}����������Dz��2�_^[��]ËU��M��B���_����;�~D�D$��+Ӄ|$ ��tM��҉T$@�l$�ۋ�t� ���Ƀ����X�u�D$@�|$ u��������t����Ƀ����Z�u�} ���  �ۍ�����������\$@���֋�t#������Ƀ����@��X����D���\��u݃}��  �\$@��+ǅ��I�������\$8��O���\$@�؋����\$(�  ���X+�����\$0����ʉ\$��	�Ã��Ƀ��D$8�������@��X����D$@�����������D���\���L$0�D$(�����D���\���\$��u����؋U�؃���  ��    +��I��ƉD$�   ;Љu�D$@��  �X�3�;Ɖt$��  �D$�t$(3�9t$�t$8�h  �D$�T$�L$(�QV�����\$P�D$3ۃ�����;��  �t$ �t$+�+�D$$�t$0����R�����I �D$$PS�u����L$P�L$(�A���M�+U�����ǃ��F�����+���+�D$3�����|Z�L$�U����������4�    ��� �Ƀ� ���A��Y��F����A��Y��F����A��Y��F����A��Y�uʋt$0�};�}"�M�� �L$�Ƀ���;��D���\��|�   ��D$ )D$$�+�;\$�t$0�����t$8�l$��;t$�t$8������M�D$@�   )\$)\$(��    T$�T$�;ЉT$�c����U�;D$@�<����_^[��]�����_^�[��]����������������U������   �MS�]�C�U,����CV��W���������������T$P�A�K��	���A�K���T$�A��A�����������������T$@��t��E0��t��E4��t��E8��t��u<�}@�V�V��W�W�������������������Dz������3�_^[��]Å��������T$8�E���E ���E�����������T$(�D$@�����T$H�D$P�����T$X���������������T$0t����ɋE0��t
��$��������H'�����H<��������AuJ������4����Az*�����T$���T$ t����̋E0�̅���   ���   ��3�����_^[��]�������������Dz;������������A� ������O� �T$ �M�����T$�E�D$�������   ��������������z���������� ��$�D$0������$�����T$ ����������Au���T$ �D$(�M�����T$����������������   ����������z���T$�E�D$���������ɋE4��t����̋E8��t�������������������������'�������8  �D$83��T$���D$H�����\$`�D$@�����M �����T$8�D$P�����M�������T$H�D$X�������T$X���T$(�T$0����M����D$H�D$8�D$X�������Ʌ�t�D$��D$ �D$`��������������������u��������������������������Ʌ�����ݜ$�   ��   Q�؃���$�   �$P�5���݄$�   ��P��$�   QS���T$|�$R���������7������P�V�H�N�P�V�H�N�P�ΉV�^����T$0����������   �؃�������$�8�����T$�M�   ����   Q�؃��D$t�$P����݄$�   ��P��$�   QS����$�   �$R�g��������������P�W�H�O�P�W�H�O�P�ωW�����T$(��������z�؃�������$������T$�M�	�T$�M�ك����T$�7���3��؉D$�D$�E(P���g������5����u�D$   �M(Q���E������5�����   t�D$�|$ ud��u*W���������5�����/  �D$(�\$0����At:�E(VP�L$pQ�I������H�O�P�W�H�O�P�W�@�G��   ��uG�U(R�D$lWP�������P�V�H�N�P�V�H�N�P�΃��V�����   _^[��]ËM��������D$@�\$P����Az!���S�V�C�F�K�N�S�V�C����A�F�Q�V�A�F�Q�V�A�ΉF�C����M(VQ�T$pR�d������P�W�H�O�P�W�H�O�P�W�σ�����_^�   [��]�������������U���,�  3ŉE��U���SVWt��} �]u	�E��M���d  �E���X  �} �Ku��9M�D  �u���9  ���1  ��]��������   輶 3�9}�e�}���  ������������Dz%hX���h@���h{  h(��.�������  ��   9E��E��Z  �U��    �E��	�����E��ɋ�u��މM�~��������D�  ��3�����E��U�|q�Q�ǋ��K���+�����    �]��B�� �˃� ���@����������D����@����������B����@����������B����@���������u��M�]�E�;�}$�ы�+�+M�����������@���������u�����詊 �E��M��с�  ��U�yJ�ʀBu�E�U�����E����U�����Ƀ�;M�M�������}����*  hX���h@���h�  ��h(�軨�����b  �   9E�E���   �E��    �M���I �����u�3����E�|]��+׉U�S�������    �]��]�N�G�A�� �`؃� �������D��`������A��`������A��`�����ű]�E�;�}�֋�+�+M���������`�����u��y� �E��M��с�  ��U�yJ�ʀBu�E�U�����E��U���;M�M��,����}�������E�3҃�|*�E�O���������    �@��� ���@��@��@�u�;�}�E��Ѓ�;�|��E���e�_^[�M�3��Q� ��]���2��e�_^[�M�3��9� ��]�������������D$�D$������z��������������̋D$�L$�A�T$,�H� �	���A�L$�H���A�H� �	���A�L$�H���A�H� �	���A�L$0�HQ�L$,R�T$,��Q�L$,R�T$,Q�L$RP�D$$���\$�\$�$PQ�������<����̋L$�D$�D��L$���D���������Dz���������������������������4��4������Au���������������̋D$�L$�D����̋D$�L$V�t$3҅�W�|��  �L$���  ;���   ��|H�T����$    �B�Z����DzX��Z����Dz?�B������Dz8�B��Z�����Dz0���� ��Å�~$�D��������Dz��������������+��G����4κ   |E�N��    �A������Dz_�A������Dz@������Dz=�A�����Dz9���G��� ;�|�;�}+�������Dz��;�|�_��^Ã�_��^Ã�_��^Ã�_��^�U�l$��u)9l$u9l$th��h��jh|�赤����3�]ËL$S�\$�����W+�3���|]��+у���V���t�����F��^�����z���F������z����^����z���F�^����z���� ��u�^;�}��I �D���\� ����z����;�|��_[]��SU�l$����   �\$����   �D$�D��VW��|$�p���+ƃ��   |z+�������T��4��d$ �B��Z�����z
�B����\���B������z	����\����Z����z
�B���\���B�Z����z
�B���\���� ��u��|$;�}*��$    �D���\� ����z�D� ���\����;t$|�_^��]��[Ã|$ u�|$ u]�[�h��h܏h�   h|��������]2�[��������������̋D$�D$�L$SU�l$ V�t$(W�|$+������\����   �W�;�}��|A�L���A�Y����DzX�A�����Dz?��Y�����Dz8�A��Y�����Dz0���� ��Å�~7���\������Dz������ ����������~������z%�~3����$WS�����ȃ���}$_3ɍ1^][Å�}��������Dz����+��ƍG�;�|�O�_�1^][Å���   ���D$ |>�T���B������Dzl�B������DzC�������DzE�B�������DzF���� ��ƅ�~:��������Dz.�����_�؍1^][�_�؃��1^][�_�؃��1^][Ã���_�1^][��������̋L$��SVW|E�t$�\$+�;�7�|$��t/;�}%��T���d$ ����;�}���\������D{�_^��[�_^���[����������V�t$����   �T$;���   �L$����   ����   ���F;�}2�^ÍD6�;���   �D���d������4���D���d������������Au�����+֍t6����T�t"�A���!��b��������At������u��ذ^���2�^�hH�h0�hq  h|�������2�^�������������V�t$��W~W�|$;�|O�T$��tG�L$��w>��S�t��u�D�������D{2ۃ�t��u��D���\������D{2ۊ�[_^�_2�^����������S�\$UV�t$�l���}^]2�[�W�|$WSV��������|9��|4;�|0���N���;�u#�D�������Dz�D���\������Dz_^]�[�_^]2�[��U����j�h��d�    P��hSVW�  3�P�D$xd�    �u����  �];��w  �}���l  �E�E���������U  ���$���������A  �E���$�ɪ�������(  �D���\������A�  �D�����$蜪��������   �D�����$肪��������   �D�����\$�L$D�D���$�|����E���\$�L$4�EǄ$�       �$�X����D$$P�L$8Ƅ$�   ������t9�\�3���~/�d$ �����L$<�$螪�����L$,�$�O�������;�|ՍL$$�Ƅ$�    ������L$4Ǆ$�   ����������ËL$xd�    Y_^[��]�h��h��h(  ���ht�h��h"  h|��M�����2��L$xd�    Y_^[��]�����̋T$��V|0�t$;�|(�D$��t �L$��t�D����L$��t�D����^�2�^��̋D$��V|:�t$;�|2�T$��t*�D0�3Ʌ�|�ʃ���;����\�����\�~�^�2�^���������U������4�ESV��W�}��������\$7�D$8},��tWh��P�y?������t	2�_^[��]��d���_^[��]ËM;�}!��tWQh|�P�E?������t�2�_^[��]Ëu��u��th\�P�?������t�2�_^[��]ÍD�3ۅ�~+��I �ރ��$��������tl�E���D�;�|݋M�D���\���\���W��\$<����Atu�D$8��t%����$�O���Q���$RWh��P�>����$�|$7 ����2�_^[��]ËD$8��t�ރ��$Sh̑P�b>�����|$7 �����2�_^[��]��D���Q�������At+�D$8��t��D�����$�y���W���$RQh`��s����E�L��ɋ֍^t��������Az7������u�M����T$<t��������zQ������u�_^�[��]ËD$8�������+��M���$���O�Q���$���Wh �P�=���� ������\$8��������E����$+���P�R���$���PWh�S����������̋L$2�����   �T$����   W�|$;���   SU�l$��Vt��uX�B�3ۃ�|7�p������Q��    ���� ���Z����Z����Z����Z�u��T$;�}�I ����;��\��|���t��ug�\:��׋�+�|;��+�������D����I �D���� ���X��D���X��D���X��D���X�u�;�}���    �D����;��\��|�^][_����������̋D$��VW��   �|$;���   �t$����   �ȃ���   ��t)�L �;�}Gh��h��hV  h|��Ș����_2�^Ã�}!hH�h��hP  h|�袘����_2�^ÍH�S�΍\�������t��+��I ���@� �@�D��u�ɋ�t��+�����D��$�@��@�u�[_�^Ã�}!h�h��hG  h|��(�����_2�^�_�^�hܒh��h@  h|�������_2�^�����������SV�t$2ۃ�|U�L$;�|M�T$��tE���D$������Au2�F�;�|������Ƀ�;��T����|���j��RQV�j�����^�[�����^��[����������V�t$2����h  S�\$���Y  �L$;��M  �T$$��U�l$ Wt	����   ��t'�D���D$ �L$���\$���$jVUPSQ��%  ��(�C�3���|;�P������N�<�    ���    �ƃ� ���Y����Y����Y����Y�u�;�}�ƃ�;��\��|�T$,�L$���t	����   +˅���4�t.�L$ �D�������\$���$j�V�T� �D$,RQSP�@%  ��(�|��C���+ȃ�|=��+Ѓ��������ۍL���<���I �ƃ� ���Y0���Y(���Y ���Yu�;�~�ƃ�;��\��_][^��������QU�l$����  �L$����  �D���D$����������  �T��������  V�t$��t/��|9\$}$h0���h�h�  h|�萕����^2�]Y�W�}���������|$�P���t����������u����6  ��    P���ˋ��ō�R��Q��} �T$,�D$$�D$0�L$(���d���t���<�������ٍ�    +Í��D$����+Ջl$ ����ul����   �D$������D$��D$��+��&+�����&��������������t�B�����������������u������u�_��^�ذ]YÅ�t[�D$������D$��D$�+���+�����&��������������t�B�����������������u������u�����_^�]Y���h�h�h�  h|��������2�]Y����̋L$����SU�  �\$4;��  �l$@����  �D$,V�t$@��t0��|9D$<}%hD�h4�h�  h|�蕓����^]3�[���W�|$0;�|&h��h4�h�  h|��g�����_^]3�[��ËD$L��t� �3��D$(Pj���$U��SP�U��������l� �D$�l$Ht���L$@�ΉT$D+\$�T$8j USR�\$L�~����L$ ����u:�D���D$(��������z+�D����������uh����h4���h  �H����D$(��+�;ȉD$u2�T������Au'�D����������Azh|���h4���h  �����D���r��D� ��$������u���d� ��������Az
�����D� ����d������������Az
���D���T$(�D� ����S�3ɉT$����Dzv��|@�T���R����D��   �R����DzK�����DzG�R�����D��   ���G��� ;�|�;���   +�t� �����D��   ����;�|��~���y���t�D��������Dzg��|@�t� �����DzU�V����Dz͍
�T�����Dzč
�T�����Dz,���G��� ;�|�;�}эT� �����Dz����;�|����+��؋L$L�ɋǉD$t�T$Љ��������L$8�\$��T$4������R�_O��������uh\�h4�h>  �Q����D$��PUW3��ay ��9t$DtR�L$ك|$8 �4�~B�T$8�\$D��T$�D$4���PSU�(y �D$L���؋D$@������l$ű\$43��D$(�D$8���$WVSP�9�������t�l$��t�L$@�4΃����|$ ŋ��ڍ׋��|$@���م�Ήl$�D$�T$ �  �D$8�l$<�T$�t$�L(�х�t'��؋�+Ë\$H���Ӎ�����Z����u���\$H�D$�L$��L$���R��R��P�4x ���|$D ��   �E��D$@���t7�l$@�\$D��<��ÍI �D$4���PSW����w ��+�+݅�u��L$�T$8�,��~7�t$4�D$@�|$D�\$ ���    ��L$8�VSW�w |$D��ރ�u�T$R�M���D$��_^][���hD�h4�h�  h|�踎����]3�[���������������̃|$ U�l$VWt���D$�L$�T$ ��S�4ʋ���    ��    P��+�QV+��w ��    �D$(�|$(��������+���������+Ã�[u��_��^�ذ��]����˅������������������t����Ƀ��@���������^u���+�+��؃�u���_��^�ذ��]���̃���T$S���\$$��UV�t$$W���t$��D�{  �l$,�����t$(�*  �ҋ�t�T��������D�  ��u����   �K�D��D$0   3��L$�D$�t$��3���|S�D$(�D$�D$0��������4�    �@��� �ʃ� �����Y��@������Y��@������Y��@������Y�u����؋D$$��;�}7�D$(�7�D$0�7ōˍËD$$��+�����ʃ������Z�u����؋L$�T$$��    D$ȸ   D$0�)D$�L$�3����t$(������D�����;t$��}A�_��^]2�[��ËT$$�t$(SUVjR�����D$<����;D$�D$(|�_^]�[�����_^]�[���U������4  �  3ĉ�$0  �} �E�MS�D$�E<VW�D$4�D$$    t��9M�L$}�M�},�O�M8���Qj P�\p �E�t$ �M�������3�;�~9]�A�t��+��\$��E,�3���=   w�|$8�P��I���M���D$$���ۉ|$t��    R��j P��o �M���E0�����E��������D�E$��   ������$������u��������D��   �D$���U�ɍЉT$��tD�\$��������ۋM�D$���+�SPV���D$�qs ����u��E�E$�E0�����������������T$(���������������������   ��~W�\$�ڋE�؋U�؋|$�ۍ�    ۉL$ �T$��I SWV��r |$,���l$u��E�|$�E$�E0�������E���E������L$�؍��T$�T$(����������������������\$��������D{C�E�����t9���D$�؋�t'���ۋ�t� ���˃�����������X�u��uك�uǃ} �܋|$���  �M��������DzG�E��W��SPQ��������u(�D$$��t	P�H����2�_^[��$0  3��;i ��]��D$(���ɋE,��t{;E�E�u�|$}�p���˃��ωT$tN��    ��+��D$ ����D$�T$ ��t*���ʃ��ۋ�t�@����b����������u��u��؃�u��|$�؉|$�}�����  �E�t$3Ƀ��D$ �L$��   �T$�J+։T$�S�������    �\$؉L$(�\$ �\$(�|��N��I �G��Y�����Dz�A��[��G������Dz	��D$���Y����Dz�A�[��G�Y����Dz�A��� �� �� ��u��\$�|$�L$;�}D�΋L$ �ΉD$��+Ƌ�+L$�D$�   �D$� �����Dz	��D$�t$փ�u݃} t�M,�UWSQR�]������}, |P�E�U8�u,��    �L$(��    �\$4��    �D$ �L$���I �T$(RWS��o \$,|$(����u�D$$��t	P��E������$<  _^[3̰�
g ��]�������������U�������  SV�uW�~�����=�  �|$$�D$@    w
�L$P�L$(�P�CE�����D$@�D$(�ȋU�����[����D$����Dz#�M�������Pj Q�%k ���_^[��]ËE������T����]����T���\$<3ۅ��\$�  �|$�E��    �����D$D����؉t$H��+��t$�|$L�|$L����+L$H�D$8�����+D$D�T$ЍA�L$<�!���L$<�M����A��M��3ɉU�D$ �7�{������   �\$�|$8�D$��|$,�}+|$���|$4�|$ �������\$�|$0�F�|$�ϋ|$,������ �� �� �x������������Z����F(�D��|$4�����x������������\��|$0���F �D��|$�����x������������Z����F�D���{�;������x������������Z����a����U�D$ �t$;ˋ|$$|�D$�t$(�<ȋ�+��D$0�Ƌt$�D$�D$8ƉD$,��+D$�D$4�D$0��ȋt$��t$,�>�t$4���l$�����������������\7���uˋt$�D$ �|$$���ʃ�;߉\$�t$�,�������4�������   ���������D�5  �xD�����A�"  ���   ��|M�r���  �V�����D��   �V�����D��   �����D��   �V����D{3ۃ��G��� ;�~�;�����   ������D{3ۃ�;�~������   ��   ��������   ��������D{�xD������Auo3Ƀ��   |=�r��t\�V�����DzR�V�����DzH�����Dz?�V����D{3ۃ��G��� ;�|�;�}��t������D{3ۃ�;�|����t������؋D$@��t	P�A����_^�[��]���U�������  �MS�]V�s��t$L�������������؍q�D$@3���   ���  W�D$Lw�|$X�Q��@�����D$L����ߍ�3�9u�L$(�ى
�t$��   �D$P��    �D$ �L$8�]�Ã��]�\$ ȃ��D$$    |X�4���������\$0ۃ�ۉ\$$�\$0��� �`��� �� �����^��A��`����^��A��`����^��A��`����^�uǋ\$$;\$ }0�t$�4��4މt$0�t$ +�\$0����`����������[�u�t$�L$8���l$ ��D�����;u�t$�L$8�#����]�D$L�u��    ���ۉT$<�u�D$$    �  �L$D���    �D$T�D$ �����D$8   ��ɸ   ��9E��D$��  �L$8�\$P�\��\$H�\$ �L$@�K�L$0�L$$����L$,�\$D�L$@����!���؋\$D��L$(���L$ �L1�   9D$H�j  �\$H+ك�����   ���\$,�T$(�D$ٍD��D$�D$$��Ƌt$�t��t$�t$(+��t$4�t$H+���T����T$���T����B��\$�b��� �� �K��\$�S�\$�H��D$ ���B��b���\$4�T��\$�H����B��b���\$�S��\$�H��D$ ���B��b��K�\$�D$ ����H���u��u�T$<�D$;L$H�	  ���ω\$�\$$ٍމ\$�\$,ٍډT$�T$(+׉T$4�T$H+ыL$����\$�a��D$����\$4�T��\$��D$����uӋT$<�  ��+ك���   �4��\$,ٍt��]�t$�t$$�T$(�4�\$,�t$�t$<�4�ٍt��\$$�t$�t$(+��t$4�t$@+�t��T����T$���T����B��\$�b��� �K��\$�S�\$��\$�D$ ���B��b���\$4�T��\$�K�\$���B��b���\$�S��\$�K�\$�D$ ���B��b��K�\$�D$ ��\$�K�D$ �����o����T$<�u;�}g���ω\$�\$$ٍމ\$�\$,ٍډT$�T$(+׉T$4��+ыL$��\$�a��D$����\$4�T��\$��D$����uӋT$<���\$ �D�L$(�L�������L$0�1���L$ �]�\1�D$@�l$D�l$,�D$0��    ��;E�ϋ|$(�u�L$(�D$������D$$t$T�l$8�D$ ��;Éu�D$$�����D$L���D$P�U����t"���ۋ�t����ʃ����^�u������uޅ�������t	P�;����_^�[��]�����������U������4  �MSVW���]�U���E�u(�D$0������+��=   �T$8�D$<    w�D$@�P��:���T$<�M���D$<�҉D$,~P�E���Ѕ҉D$4�T$(t1�l$(��    Pj V��` �E$�������|$( u֋M�D$4�E$�؍4���M���M$���Qj V�` �M��9M|�Q��U�D$,�E�UP���$RQ������M����t!�D$,�UPQ�MQR������M������   �D$0��    �A�T$4�D$(3�9U��   �L$8��    �D$0�L$,��3Ƀ�|F�C�������    ��� �Ƀ� ���F��^��G����F��^��G����F��^��G����F��^�u�;�}��+�����Ƀ����F��^�u�|$0�؍�    ��+�;U�t����M�E$+|$4�����E���D$,�l$(�0����}��   ���M$�ٍ΋u3����U(��   �B+׉T$4�S��]���D$0����    �D$(Ë\$0�t��O�D$8�F��Y�����Dz�A��[��F������Dz	��D$4���Y����Dz�A�[��F�Y����Dz�A��� �� �� ��u��U(�]�D$(�t$8;�}'+׍Ǎ4�+؋�������Dz��������u�D$<��t	P�8����_^�[��]�����������́�  SU��$0  V��$   �]���������=   W�D$    w�|$ �P��7�����D$��݄$<  ��$0  ��$,  ��$(  WV���$UP��$L  QRV�^�����$���D$to��$$  WVUP����������D$tT��|P��$$  ��$D  ���    ��    �T$�D$��$H  UWV�{a t$$|$(������$H  uڋD$��_^][t	P�b7�����D$��  ����̋T$�L$�D�������Dz]�����D��\������DzI�D$,�D$ P�D$,P�D$$���$P�D���D$(���\$�D���T$<�$R�T$,PQ�L$8QR������8ËD$,�D$ P�D$,P�D$$���|$ �$Pt�D$,P�D$,PRQ�L$(Q�8�����(ËD$(P�D$0RQ�L$$Q�������$������������U�����M,��t  SV�u;�W|	�F��D$P��L$P�];�|	�S��T$`��L$`�} �}t���E$����+ǉD$\�A��������    �L$t�ȉD$l�3��=   �|$d�D$|    �L$Xw��$�   �L$@�P�5�����D$|�D$@�T$@�D$X�4�P��j S�t$T�\$|�[ �E0�L$L�]�U��Q���$SR������E8�E��V�u���$VP�������|$P t+�L$@�T$P�EQRSP������L$X�T$p�EQRVP������ �M�ɋD$p��   �T$@�T$4�U ��҉T$X�U(�T$8�L$D���    �T$83�9]~I�4�    ���L$H�ًL$4�	��t����Ƀ������@��X�u�L$\����Ƀ�+��;]|��T$XT$8�D$4�l$Du��}, �  ��    ��} ��   �T$@�M�T$<�ʉT$4�U(�T$8�L$D�L$83�9]��   �u�����T$L�T$H�4���T$H�ڋT$4�
��t����Ƀ������@��X�u��    ��+ʅ��T$<����t����Ƀ������@��X�u�T$\��+D$L��҃�ʃ�;]|��M ���L$8�   L$4L$<�l$D�B����},�&  �T$`������L$L�L$Pу��V  �U���D$<    �C  �L$@�u�щL$T�M(�L$4�L$43ۅ���   �T$H��T$8�|$P~E���t$<�U�V�t$@�֋T$H�ڋ�t����Ƀ������@��X�u�u�؍�    +��	��    ��T$8��T$T�
��t����Ƀ������@��X�u��    ��+ʃ|$`~B���s�t$H�֋T$@�t$<���t����Ƀ������@��X�u�u�؍�    +�+U$+D$L�D$8��҃��;������U�M �D$<�D$T���L$49T$<������},��  �   9u,�t$D��  ���҉T$X�L$`�;�L$8�t$8�} �D$<    �H  �M(�L$\�} �T$\�T$4�D$h    �  �d$ �\$83�;t$P��~;���   �4�    ��ƃ�;L$P�;���   �]��L$<��\$@�ˋ\$H�L$T���ML$h�ލˉL$L�L$8�+�����х��\$L��\$T���t'���\$x�\$4����ɉ\$4�\$x�����@��X�u�t$T�����)|$4�}���|$L���|$du��M$�׋t$D���L$4�L$h����;M�ЉL$h�����M �T$<���L$\��;U�T$<������T$X����    �;u,�t$D�T$X�w����} t�T$p�E,�MRWPQ�G������l$t�\$l��~F�U@�uD��    �|$p��    �D$l�L$x��$    �T$tRWV�Z t$x�$�   ����u�D$|��t	P�0����_^�[��]��������U�������   �E+ES�]VW�D$(�E�{���    �4�F��F��T$�D$��L$0�T$ �D$,    ��������Dz)h����h����h�  hd��p����2�_^[��]Ã} �M  ���E(��������Dz$�u�����D0���������Dz�ذ��_^[��]��پ����9uu���E ��E� ������Dzs�u��9u�  ���؋T$��t�����"�������Y�u�U�؍�    +ȋE�؋����ډ]�t$��  �������+Ѝ�    �T$�D$ �2���E����~���R���H.���E(���D$�D$,���g����]�T$���|$�Ét$tY�\$(��ۋt$ �>�u�'�l$�����y�+�+Å�����t�B�������� ���������u�|$ ����u��t$�D$ +ȃ������t$�D$ �v����   �E��M�؅��ى]�|$��  ���    �D$��+ʍ4��L$�t$��]���Ë�tO�|$(�����U�����+���+ǅ�����t�A�������� ���������u������uËL$�|$�t$�������|$�t$u������؋D$,��t	P�%-�����_^[��]����E(��������Dz�E� ��������Dz_��^�ذ[��]��ڃ}u���E �D�]�����D�������Dz	�E   �&���E   ~��R���i,���E(���D$ �D$,�ȃ}��   ���؋֋�t�����������Y�u��    �؋�+ȅ҉T$�%����E��}�ǉD$ ��    +��D$�t$�D$�ҋE�|$ �t$��tT�T$�2�U�&���������y�����t� ���ʃ�����������X�u�T$(�����������u��T$�D$�   )t$t$+ȃ�+ƅ҉T$�D$�s����m����������_����E��M����    +��T$ �t$���E�T$ ��tO�L$(��ɉL$���M�&������������t� ���ʃ�����������X�u�L$�����х�u��t$�������t$u�������������U������,  �} SVW��   �} ��   �]����   �E9E��   �}�� �L$8�w��L$�D$,    ~��    Q�^*�����D$,�D$�Ⱥ   �;�~�����d��������{D��;�|����D���G��d����4����{%�U���F  �E �]��+؉t$$�\$0�T$(���2�_^[��]���I �\$0�33ۃ�|J�U�ҍw���҃�����    ��    � ��Y��� � ��Y�� ��Y�� ��Y�u܋L$;�}�U���� ���\���;�|�   ;��D$�  �]�u�O��S�L$�T$ ��$    �|$�ȉL$��   �D$�L$ �W��T��\$+������������\$��$    �B��� �aЃ� ��� ���a����H��B��&�����H����X��B��a��B��&���H���a������H����X��B��a��B��&���H���a������H����X��B��a���a����H��B��&�����H����X��j����D$�}�]�L$;�}\��+ЋD$�ЍT:��ӉT$4��+T$�L���\$4�d$ ����a���������a�����C��&�����H����X�uӋD$�]�l$�D$ ����;ǉD$������L$�t$$�����l$(�t$$������D$,��t	P��'����_^�[��]����������D$S�\$�D$U�l$V�t$ W�|$ ���\$���$jVWSUP�����D$X�L$<�\$ �D$P���$j�VWSUQ������(_^][���VW���W|���~���M|������~������~��_��^����������̃|$ ��~��� �VW��~W�c~����t���؅����t���ͅ����t_�   ^�_3�^������������̍AP�g����������V�t$QV����}����^� �����������V�t$QV���}�����������^� �������D$���A(�Y����Dz�A��A(���A�����A �Y���A��D{	�����I ���A�����Dz�������A�����������V�ʋt$���\$���\$�$��{����^� �����������̃���QS�YU�i�l$�iV�qW�y�)�i�i�i �i�i$�i�i(�i�i,�A�D$$�Q�q �y$_^�i�Y(]�A,[�����̃�@S�\$L2���V����   UV�D$ �nP���z|���L$������T$������������   W�؋|$TV���ݑ���\$U���ё���\$����u+�L$ QV�T$@R���$|�����M|���t$_]^��[��@� �D$ PU�L$@Q����{�����"|���t$_]^���$�[��@� �2�]^[��@� ������������̃�VW��L$�D$PQ�������D$�|$���$W��������_^��� �������̃� V��D$P�L$,Q��������D$���T$�$R��������D$P�L$,�Ր��^�� � �������������̃�VW�|$$��V�D$P���������P�V�H�N�P�V�H�N�P�V��V�D$P��������P�V�H�N�P�V�H�N�P_�V�^��� ���������̃�LSV��V�D$@P�N�z���D$<���D$\�L$\�����ل�t�D$\ �D$D�L$
��������A{�D$
 �D$L��������Az���2ۈL$�L$�Bx���L$$�9x���ۊL$\��   ��t�D$
��u}������� ��L$���T$���D$���L$���T$���D$ ���L$$���T$(� ��D$,�$��L$0�T$4�D$8��  �D$
����   ��t��uy�������L$���T$� ��D$�$��L$�(��T$�,��D$ �0��L$$�4��T$(�8��D$,�<��L$0�T$4�D$8�4  ����   ��t��uy�(��,��0��L$�4��T$�8��D$�<��L$����T$����D$ � ��L$$���T$(���D$,���L$0�T$4�D$8�   �D$<�L$�\$�D$D�\$�D$L�\$��}���L$Q�L$(�Cs���|$\ tu�|$
 tn��tj�L$�D$ �����tX��������\$��� ��\$�T$$�����D$(�\$� ��L$,�$��T$0�D$4�L$8�L$X�T$$R�D$PV��M���D$^[��L� ������̋D$V����P�V�H�N�P�V�H�N�P�D$�V��N�PW�~�W�H�O�P�W�H�O�PW�ΉW�w����t ���)����t�������t
_�   ^� _3�^� ���������j�h��d�    PQV�  3�P�D$d�    ��t$��  �H+���\$���   ���D$$    �$莂����ݞ�   �ƋL$d�    Y^�������H+SV�t$W�ك��\$�"   �����$���   �A��_^��[� ��������̃��D$��V�\$W�|$W��L$PQ���  ��t?��T$Rݞ�   W���4  �D$ݖ�   ����;������t��7����t��_^��� ��_2�^��� ������j�h�d�    PQV�  3�P�D$d�    ��t$���   �D$    �e������D$�����  �L$d�    Y^��������VW��j ���   �ol���|$���$W���  ��_^� ������VW��j���   �?l���|$���$W����  ��_^� �����̃�V���   j���l���\$j ��� l���l$^����������Q�D$���   ����   �P���   ���   �P�$    �HY� �������������j�hH�d�    PSV�  3�P�D$d�    ��3ۍL$�\$�l����t@�L$�0l���ؕ����z*�D$�L$ �T$$���   �D$(���   ���   ����   �L$�D$���������ËL$d�    Y^[��� ��j�hx�d�    P��SVW�  3�P�D$d�    ��3�S�L$,�\$$��j��j�L$,���j��� �����A��   j�L$,�j��S�L$,���j���� �H6����AzZ�D$(�L$,�T$0���   ��D$4�N�V�ΉF�,k���H+����Au#S���Gj��� �H+j���\$�2j���D$���L$(�D$ ���������ËL$d�    Y_^[��� ��j�h��d�    P��SV�  3�P�D$d�    �����   ��҅�u�D$,��|v��
q��Ph�L$Q����j���D$(    �i��� �\$0����Az�2ۍL$�D$$�����J�����t2��L$d�    Y^[���8 ��L$d�    Y^[���8 �ËL$d�    Y^[���8 ���̃�VW�����   ��l���D$�w0P���?u�����P�V�H�N�P�V�H�N�P�V�D$�wHP���u�����P�V�H�N�P�V�H�N�P�ωV�C��_�^���������������̃�V��W���   j���h���\$j ���h���l$_܎�   ^���������������U������SVW��M�D$PQ���b  �؄���   �ƈ   j ���9h���l$�T$�������H+��At���������������{����T$��������Az��������A{����\$����؋��h�����D$������z�����T$������Au'����$��$������z���\$����\$������؋}��tj ���g���D$�_^��[��]� ��VW����  ��tT���   ���Si����tCj���Fg���\$j ���9g���l$��;����Au�������H6����Az_�^���_2�^�������j�h��d�    P��  UVW�  3�P��$�  d�    ���D$    ��$�   �   ����m���� ��y�L$������$�   �T$�D$@�L$<R��Ǆ$�     �D$4�������$�  Vt�L$�g�������  �L$�D$   Ƅ$�   �5����Ƌ�$�  d�    Y_^]�Ĭ  � �������̃�V���   j���f���\$j ��� f���l$^���%H+����;����Az����2��������������V�D$W�ы����   ������z����T$�����$�pw�����Y�����ݟ�   ���Hf�����H+_^����Az�� 2�� �������������j�h(�d�    PSUVW�  3�P�D$d�    ��t$$�    �����D$    ��\?���D$$�L$(݀�   �T$,�D$0ݝ�   ���   ��L$4�V�F�N���Df����t��2���h�����������e���H+��������z�2�ݝ�   �����t	���/����؍L$(�D$�����L����ËL$d�    Y_^][��� ����j�hf�d�    P��   SVW�  3�P��$�   d�    ��݄$�   ���\$�L$ ���$��x����݄$�   ��$�   ���$P�L$,Ǆ$�       ��  ����̉�V�Q�V�Q�V�QP��Ƅ$�   �p����L$ ��Ƅ$�    �  �L$Ǆ$�   �����i����Ë�$�   d�    Y_^[�Ĥ   � ������������U����j�h��d�    P���   SVW�  3�P��$�   d�    �ى\$ �L$<�  ��u�\$$�E�MVPQ�L$HǄ$      �	  ����   �T$$RV�L$D�  ��to���D$$������Aud���\$�L$<�$�w������̉�P�Q�P�@�Q�A�L$LQ��Ƅ$  �M������L$,��Ƅ$    �W�����ta�\$ ����ع    ��Z���ݓ�   �����   �T$�$�0t���L$<Ǆ$   �����L  2���$�   d�    Y_^[��]� �L$<Ǆ$   �����  ���$�   d�    Y_^[��]� ����j�h��d�    PQV�  3�P�D$d�    ��t$�D$    �  �H+���\$���   ���D$$�$�yv���L$ �T$$���ĉ�L$8�P�T$<�H�P�D$,P���D$(�����L$ �D$�����'����ƋL$d�    Y^��� ��j�h�d�    P��SV�  3�P�D$d�    ���D$0���\$�L$���$��u������̉�P�Q�P�@�Q�A�L$<Q���D$8    �����L$���D$$����莯���ËL$d�    Y^[��� ��������j�hV�d�    PQV�  3�P�D$d�    ��t$�c   �H+���\$���   ���D$$    �$�.u���D$ �D$���$P���D$ ������ƋL$d�    Y^��� ��������������V���(9����ݞ�   ��^�������������黮�������������݁�   ���������̍AH�������������U����j�h��d�    P���   SVW�  3�P��$�   d�    �ٹ    ��|$d�uV��Ǆ$�       ��?�����D$u�    �t$d����  �D$|P�L$8Q��������{W�L$8�h���\$�C0P�L$8�h���T$�D$����������������A�0'�H<z\�����T$$����������   ��������z���T$����\$�����T$��������Az|���\$����������Azw�\$$�s�����T$$����������z���T$����\$�����T$��������Az5���\$����������������Az"�\$$����������������������������؍�$�   R�D$PP��������L$4�P�T$8�H�L$<�P�T$@�H�L$D�PW�L$8�T$L�Cg���\$,�C0P�L$8�2g�������D$,����������Azd�����������  ����������z����0'���������H<����������   ������������������A��   �����Y��������������z����0'���������H<����������   ������������������Azv�������������D$������Dze��������DzZ���D$$�����T$,����������4��������   ������������D{I���D$,��$�;��������������������D$$�����L$���L$�����������{1 ������������Au)��$������4����Au܋�   ݛ�   �����؍L$dǄ$�   ���������D$��$�   d�    Y_^[��]� �j�h��d�    P��  SUVW�  3�P��$�  d�    ��L$\��b���L$��b���L$,��b���L$D��b����$�  ��$�  ��$�  SVW�L$P�|z������  �D$DPW��$  �R:��V��$(  Q��Ǆ$�      �d��PV��$t  R���Fd����$P����$  �$P��d����P��$�  ��9��V��$X  Q��Ƅ$�  �4d��PV��$�  R����c����$P����$L  �$P�d����P��$�   �9���L$\Q��$�   R��$�  P��$  QƄ$�  �O�  ������   �T$\R�D$xP���c����L$�P�T$�H�L$�P�T$ �H�L$$�P�L$�T$(�h��ݕ�   ��������zZ�L$��h����tM�D$P�L$HQ�T$|R��j����L$8�P�T$<�H�L$@�P�T$D�H�L$H�P���L$,�T$@�zh����u\��$�   Ƅ$�  袨����$�  Ƅ$�   莨����$  Ǆ$�  �����w�����    ��Z���ݝ�   2���   �D$\�L$`�T$d�E �D$h�M�L$l�U�T$p�E�D$�M�L$�E�D$ �M�L$$�U�T$�U �T$(�E$�D$,�M(�L$0�E0�D$8�M4�L$<�U,�T$4�U8�T$@�E<�D$D�M@�L$H�EH�D$P�ML�L$T�UD�T$L�UP�T$X�ET�MX�͉U\�+3����$�   Ƅ$�  藧����$�  Ƅ$�   胧����$  Ǆ$�  �����l������$�  d�    Y_^][�Ĕ  � ��������������V��݆�   ���$�X������t��ܞ�   ����z���_5����t�^�2�^�����D$VW����E ܎�   ���$�D$�D ܎�   �|$���$W���1����_^� ��������������̃�SV�t$ ��W���   �D$P�T$R�T$(�:���ĉ8�z�x�z�x�z�x�z�R�x�P�b2���������D$��������D�D$z��������Dz�ي����_^[��� ��� V �����������Au�H+�_^[��� ��_^[��� ����������̋D$�D$P���$��;��� ���������j�h�d�    PQSVW�  3�P�D$d�    �ى\$��/���t$$�    �����D$    ��3����u����0���D$(��ݛ�   �L$d�    Y_^[��� ���������j�hO�d�    P��|SUVW�  3�P��$�   d�    ��3��|$��$�   �ˉ�$�   �i�����$�   �D$   �|$0�   ����I]������y�݆�   ���\$�D$(݆�   ���$P�/��݆�   ����L$0�P�T$4�H�L$8�P�T$<�H���\$�L$P�P݆�   �D$(�$P�ΉT$X�R/��݆�   ��L$H�P�T$L�H�L$P�P���\$�T$d�H݆�   �L$h���P�$�D$(P�ΉT$p�/��݆�   ����L$`�P�T$d�H�L$h�P�T$l�H����$�   �T$�P�$�D$(P�Ή�$�   �.����L$x�P�T$|�H��$�   �P��$�   �Hj ��$�   �P�D$4Pjjj j�ˉ�$�   �ͽ���Ë�$�   d�    Y_^][�Ĉ   � ���������������j�h��d�    P��d  SUVW�  3�P��$x  d�    ��L$x�D$ �[����$�   �w[����$�   �k[���L$H�b[���L$`�Y[���L$�P[����$�   �D[���L$0�;[����$  �������$H  Ǆ$�      ������$�  ��$�  W��$�   P��Ƅ$�  ��\�����$�  �L$x�P�T$|�H��$�   �P��$�   �H��$�   �PS�D$|P��$   Q��$�   �3d����T$$�H�L$(�P�T$,�H�L$0�P�T$4�@���L$�D$,��a�����m  U��$�   Q���&\����$P����$�   �$R��\�����$�   �P��$�   �H��$�   �P��$�   �H��$�   �P�D$(P��$�   ��$�   Q��$�   R�wc�����$�   �P��$�   �H��$�   �P��$�   �H��$�   �P����$�   P��$�   Q��$�   ��$�   �][��P��$�   R��$   �����D$P��$�   SQ��b�����$�   �H��$�   �P��$�   �H��$�   �P����$�   �@��$�   Q��$�   R�ω�$�   ��Z��PW��$P  �B�����$  P��$�   Q��$P  R��$$  P��  ������  ݄$�   ����$�   �$Q��$$  �!�����T$0�H�L$4�P�T$8�H�L$<�P�T$@�@�L$0Q��$�   R�ωD$L�tZ����L$H�P�T$L�H�L$P�P�T$T�H�L$X�PW�L$4�T$`��o��ݞ�   �L$H�_�����1  �D$HP�L$Q��$�   R�a����L$l�P�T$p�H�L$t�P�T$x�H�L$|�P��S�L$d�T$x�Z����$����z�L$�_���L$`��^����$�   ��^���D$0�L$4�T$8��D$<�N�L$@�V�T$D�F�D$H�N�L$L�F�D$T�N�L$X�V�T$P�V �T$\�F$�D$`�N(�L$d�F0�D$l�N4�L$p�V,�T$h�V8�T$t�F<�D$�N@�L$�FH�D$$�NL�L$(�VD�T$ �VP�T$,�FT�NX�ΉV\�$*�����]�������\$��$H  Ƅ$�   聞����$  Ǆ$�  �����j����Ë�$x  d�    Y_^][��p  � ������������U������4S�]VW3���|$ ��`�D$ �8'��$�T$ �= ܎�   ���$�D$(��; ܎�   ���D$8�$P����(���L$(�T$,���ĉ�L$H�P�T$L�H�L$P�P�T$T�H�ˉP�Kb�����]����At�����|$ �i����_^[��]� _^2�[��]� ���������V���'����ݖ�   ��ݞ�   ^�������݁�   ����݁�   ��������Az3���   ݄р   ���$��������z"�ظ   +��������������9# �$������������%# �$����������������̃�8VW���t����T$݆�   �~ܞ�   ����A{�~0W���D$�$P�W����P�L$,Q���V���D$��L$D��P�Q�P�Q�P�Q�P�Q�@W�A���L$4�$Q�KW����P�T$R���V����L$H��P�Q�P�Q�P�Q�P�Q�@_�A�^��8� �������������������������̃�VW3�Wh � @���������D$u
_3�^��� �D$=����|$��v�����T$ S+�U��@@  �荞<@  ʍF<��L$��H@  ǆL@   @  �D$$   �|$(��$    �|$$ �  ��u9�@@  u�D$(   �D$(PS�v�  �Ѓ��҉T$��   � @  +�L@  t3�F<PW����������D$��   |$�T$�F<��H@  ǆL@   @  �|$(u	����   ��vW��@@  �����sI��t"�; t����+�;�v���+�D$��@@  �,�������v�����L$+�D$���@@  �	��u�l$$���	����!h�h��h,  h���?�����D$ ���O����][t�D$�|$ u	�D$ �D$��_^�#D$��� ����̃�SUW��D$3�P�L$Q��3��\$�\$ �\$$�\$(�C����u&�L$,;�t�D$(;�vPSQ�7# ��_]2�[��� �|$ � @V�t$,u>9\$$|8�D$ ��v-;�v)9\$0t#�x�W�������;ÉD$tPW��������D$,��\$,�]4��������u�D$,9]4�\$0��#T$,��u��t��vVj S�" ���|$, u�D$��t	P������^_]2�[��� �������v�����L$��<@  �+��������@@  �L$��v�������H@  +���L@  �T$�D$0   3ۍd$ �|$0 �/  ��u9�@@  u�   ��<@  SP��  ������   ��u	����   3���vV��@@  �����sH��t9�<@  t����+�;�v��ȉ�@@  ��������v�����L$��<@  ��@@  D$+���ve��L@  �����sW��t)��H@   t ����+�;�v��D$ȉ�L@  +��#����������v�����T$D$��H@  ��L@  +��������������l$0�����hl�hL�h�  h���N<�����D$, �D$��t	P��������|$0 u�D$, �D$,^_][��� �����������V��F8�����w$�$�@p��<@  P�O�  ���<@  Q�1�  ��j8��<@  j R�n  ���F8    ^Ë�pp"p"ppp��������SVW��2��$�����tR�~8�Ä���   ���j���j8h����<@  j	W�U�  ����u_�F8   ^�[�j8j W�� ��_^��[Ë�跟����t9�~8�Ä�u5������j8��<@  h��W�^�  ����u�_�F8   ^�[Ë������_^��[��������������QV���D$ �b�����u^Y� U�l$W�|$��v��t1W���_����t%��u	_]�^Y� UWj �7����P���������u	_]2�^Y� ���   S�Äۈ\$t���������u���I���2ۈ\$�D$P���g�����u[_]^Y� �Ã� t(��u0UW���u��������D$�����D$[_]^Y� UW�������D$�D$[_]^Y� �̃��D$S2ۅ�V���D$    �\$t�     �H�����u^[��� U�l$��u]^�[��� W�|$ ��t,�D$P���������t�L$Q��������t�D$��t<t_]^2�[��� ���� t&��ul�������؄�tWU���d����؋��+����WU�������؄�t<WUj �!6����;D$t*hЖh��h�   h����8���D$4����t�    _]^��[��� �̡����$��uD�$�D$�D$�D$�D$�D$�D$�D$�D$ �$P�4!�D$�����w
�   �����$������������̋��     �@����ËT$���L$��P� �������������̋L$3���3wjtb�����(��   ���t�$��t�   ø   ø   ø   ø   ø   ø   ø   ø   ø   ø   ø)   ø3   Ã�dw;t3��Ã�wd�$��t�=   ø>   ø?   ø@   øA   øB   ød   Ã�gwt��et	��u"�Aføe   øg   Ã�ht���u�øh   ÍI �s�s�s�s�s�s�sttttt�t 	
�I ;tAtGtMtStYt�����������̋D$�T$��Q� h@jj��(Q�@B ��������������V�t$Wj j��h � @���hy����u_^� �SP��������؄�tS�OXQ��������؄�tB�WRj��������؄�t/�G(P��������؄�t�O8Q��������؄�t��HW�������؋��d����u2ۊ�[_^� ������V�t$Wjj��h � @����x����u_^� SW���&����؄�t[�GP��������؄�tJ���   Q�������؄�t6���   R��������؄�t"��(  P��������؄�tV��0  ������؋������u2ۊ�[_^� V�t$Wjj��h � @���(x����u_^� SW�������؄���   �GP�������؄���   �O Q���l����؄���   �W(R���7����؄���   �GHP���B����؄�tp���   Q���.����؄�t\�WPRj���+����؄�tI���   P��������؄�t5�OpQ���6����؄�t$���   R���"����؄�t�ǐ   W�������؋�� ����u2ۊ�[_^� ������̃�V�t$3�W�D$�D$���D$P�L$Qh � @��������u_^��� �|$S�Ä���   W�������؄���   �WR�������؄���   �G P���6����؄���   �O(Q�������؄���   �WHR�������؄�t~���   P���8����؄�tj�OPQj��������؄�tW���   R�������؄�tC�|$|<�GpP��������؄�t+���   Q�������؄�t�|$|�ǐ   W�������؋������u2ۊ�[_^��� V���   W3�;�tc���~� ��Wu9�8���   ;�t	��Pj�ҋ��   ;�t	��Pj�ҋ��   P�������hD�h�h3  h��2�������   ���   ���   �~_^�����̡`/��V���d/�N�h/W�V�l/���N�$�F������`/���   �d/���   �h/���   �l/���   ��3��$���   ���   �a���h@h`�jj��X  ��(  ǆ,  ����R��0  ��4  ��= �5���  ǆ�  ����ݖ8  ݖ@  _ݖH  ��ݞP  ^���������S�\$��U��~dW�|$��|ZV�t$��|P;�tL�E�;�B;�>�M�;�~�;�}��P���֦���Eiې  i��  i��  S��WV�U ��^_][� �����������V��~ ���t%�F��tj P����F    �F    �F    ^�����������VW�|$��;�tA�G��_�F    ��^� 9F}P�4����N��t�G�Fi��  P�GPQ�F ��_��^� ������������V��L$��|9�F;�}2+���P�APQ�������F��Fi��  Fh�  j P�� ��^� �������̋D$�L$i��  PQ�������� �����V��~ ���t%�F��tj P����F    �F    �F    �D$t	V�/�������^� �����̃�`VWh@h`�jj�D$@3�P���t$�t$ �|; �5�T$h@�T$�t$d�T$$j�\$0�D$l�����   �t$�j�L$<Q��: _^��`�̃�VW�������|$3��D$�D$�D$P�L$Qh � @����	����u_^��� �|$S�Ä�taV���O����؄�tS�VXR���~����؄�tB�FPj���;����؄�t/�N(Q���*����؄�t�V8R�������؄�t��HV�������؋��o�����u2ۊ�[_^��� �������������̡`/V���d/�N�h/�V�l/�FW3��~�~�~�F�����~ �~$����N(����V,����F0����N4���h@h`��V8���jj�Np�F<�~@Q�~H�~L��9 �5���   ǆ�   �����VP�VX���V`�^h���   ���   ���   ǆ�   �����   ���   ���   _^�����������V���h����`/��d/�N�h/�V�l/�F3��F�F�F �F$����N(����V,����N0����V4����N8����V<�F@���   ���   ���   ^�������������SU�l$��;���   VW������E ��M�K�U�S�E�C�M�K�U�S�E�C�M�K�U �S �E$�C$�M(�K(�U,�S,�E0�C0�M4�K4�U8�S8�E<���   �R�C<�M@�K@�uH�{H�   󥍋�   ���   P�ҋ��   ���   ���   ���   ���   ��_���   ^t�}  ��~�E ][� ��][� �������������j�h��d�    PQSVW�  3�P�D$d�    ���|$�D$   ����3�9��   ���   �\$���t�F;�tSP������^�^�^h@jj��pW�D$,�����7 �L$d�    Y_^[����������́�  �  3ĉ�$�  VW���L$����h@jj��$l  �d   �t$P��6 ��$�  _^3�� �Ĕ  �������̃�VW�������|$3��D$�D$�D$P�L$Qh � @�������u_^��� �|$S�Ä�tpV���/����؄�tb�VR�������؄�tQ���   P���
����؄�t=���   Q���ֺ���؄�t)�|$|"��(  R��������؄�tW��0  �	����؋�� �����u2ۊ�[_^��� �����������������V���T$���T$�N�$�    �oH������T$�T$�N0�$�WH������T$�N�$�3H���NH��t��Pj���FH    �NL��t��Pj���FL    ^����V�t$Wj j��h � @���hl����u_^� �SP��������؄���   �OQ�������؄���   �W0R�������؄���   �GP��������؄���   j jh � @����k���؄���   �H ��Q�������؄�t�H t�OH��B V�Ѕ��Ë��/�����tP��tNj jh � @���k���؄�t8�L ��Q���R����؄�t�L t�OL��B V�Ѕ��Ë��������u2ۋ��������u2ۊ�[_^� ����j�h�d�    P��SUVW�  3�P�D$0d�    ���"����t$@�D$(P�L$ Q3�h � @�Ήl$(�l$4��������  �|$�Ä���  �T$ R�Ήl$$�V����؄���  �D$ �����w5�$�ԅ�   �&�   ��   ��   ��   ��   �GP�������؄��S  �O0Q���˸���؄��>  �WR�������؄��)  �D$$P�L$Qh � @�Ήl$$�l$0����؄��  �|$�D$@ �Ã����tT�T$@R��������؄�tB�|$@ t;j,�������D$,���D$8    t	����t���3��GH��ȋB$V�l$<�Ѕ��Ë���������   ����   �L$$Q�T$Rh � @������؄�tf�D$P���D$ �X����؄�tB�|$ t;j@��������D$,���D$8   t	���S���3��GL��ȋB$V�l$<�Ѕ��Ë��)�����u2ۋ�������u2ۊËL$0d�    Y_^][��(� ����'�/�7�?�����j�h;�d�    PQV�  3�P�D$d�    ��t$�N�@2���N�D$    �p9���N0�h9�����FH    �FL    �����ƋL$d�    Y^���j�hk�d�    PQV�  3�P�D$d�    ��t$�D$    �;����N�D$����蛀���L$d�    Y^�������������VW�|$��;���   ��������O�N�W�V�G�F�O�N�W�V�G�F�O �N �W$�V$�G(�F(�O,�N,�W0�V0�G4�F4�O8�N8�W<�V<�G@�F@�OD�ND�OH��t�[T���FH�OL��t�LT���FL_��^� ��U����j�h��d�    P��  SVW�  3�P��$�  d�    ������u�]�����N����V����F����N����V�C�K������  �$������  ;O��  �I�O��R���8����  ����  ;�T  ��  ���P  �y ��  �I����  �����  ;G��  �O�@��R���=8���  �{H�y  �CX�CP�%�$����4����A�Z  Q��$�   P��8  �4����$�   Ǆ$�      �ĺ����t?�CP����$\  �$Q��$�   �3������H�N�P�V�H�N�P�V�@�F��$�   Ǆ$�  �����*~����  �{H��  �CP�CX�C`�Ch�%�$����4����A��  ����  ;O ��  ��O�ً���~  �O;��s  �C���h  ;��`  �C���U  ;��M  �C���B  ;��:  h��jj�L$@Q�L�����@�G��Q�L$8��6���C�@�G��Q�L$P�6���C�@�G��Q�L$h�6���[�G�[��Q��$�   �6���}�Gh�T$|R����$H  �$P�8���G`��P��$p  Q�T$lR����$  �$P��7���GX��P��$�   Q�T$\R����$@  �$P�7���GP��P��$�   Q�T$LR����$0  �$P�7�������6�����6�����6�����P�V�H�N�P�V�H�N�P�V���~>����$�  d�    Y_^[��]� ����h������V��F���    �F    tP�������F    �F���F    t�0P�c���������u�^���������SVW�|$��;~�~+�N���PQ�O��������Fu_�F�^2�[� �~_^��[� �������������S�\$�C�=�� V��w�;N|�	��;�}��P��������u^3�[� ��V�@U����,�    W�E�<�P��d����؃���u_]^[� �L$�CU��h�   P�G�W�X �F�����_]�^^[� ���̸�������������j�h��d�    P��VW�  3�P�D$ d�    ��t$��[���D$3�P����|$,����������N�P�V�H�N�P�V��/�F��/�N��/�V ��/�F$�F(   ���   ���   ���   �ƋL$ d�    Y_^�� ����������������V����]�����   ��t)W�>3Ʌ�~�VS�������Yu�[�V�QʍD�_^����QVW�|$j��jh � @�ωt$�Ca����u_3�^Y� ���   ��SUu3���(����   �8 ��   �p��u3�U��胿�������   ����   ���D$    ~O��I �P���V����؄�tb�N�QR���2����؄�tN�F�PQ�������؄�t:�D$����;ŉD$|��t$���   R�������؄�t���   P�������؋��������u2�]��[_^Y� 3��B�����������������̋L$hܗ������   � ���������̋��   ��t�8 ~�   �3���������̃�VW�|$��;��t$��   S�3����;^~%�N�[��PQ����������Fu�F���^3�9�D$�}   �D$U�d$ �GD$�X�ۋh�0t?��t;�L$V�o�������t'�G��    RSP�G �W������QUR�5 ���|$ �D$�D$��;�D$|��D$][_^��� [_��^��� _��^��� �������j�h��d�    PQ�  3�P�D$d�    h�   �u������D$���D$    t���k����L$d�    Y���3��L$d�    Y�����������̃�UVW�����   3�;��|$t�������V���������   �|$$�D$P�L$Qh � @�ωl$ �l$(�@�����u_^3�]��� �|$S�Ä��  �T$R�ωl$蠫��9l$���   ����   j蕿����;�t�(�h�h�h�3�;ŋt$���   ��   �L$Q���q���9l$�l$��   �I �T$(R�ωl$,�0����؄���   �D$(;�~H���   P������;�tI�F�L$(PQ�������؄�tb�V�D$(RP���֪���؄�tL�L$(��t$�D$��;D$�D$|���t$�|$ |$���   R��說���؄�t���   V��薪���؋�������u2���[_^]��� ���������̋D$V��3ɉ�N�N�N9~9HtP���������^� �����S�\$V��;�tuW���   ��t�������W�,�����ǆ�       S���W�����    _t&j��������t���   Q���q����3����   ���   ���   ���   ���   ��^[� ��������j�h+�d�    PQVW�  3�P�D$d�    ��h�   葽�����D$���D$    t���������3����D$����tW�������ƋL$d�    Y_^������������VW�|$��t5h����������t%�t$��th����������tW������_�^�_2�^�������������V��W���   �����t������W�Ͼ����ǆ�       ����U���D$t	V设����_��^� ���̃�0S�\$8U���   ���*8����t�|$@ uD���hs����聝����t2VW�D$P��������   ���L$�+s��_��^ݓ�   ݛ�   ����7����]��[��0� �������QV�񋆈   ����L$~>S�\$UW3��萋��   ��SP�Bt���Є�u�D$�Ǩ   ��uڊD$_][^Y� ��^Y� ������̃�S�\$U�k$V��NxW�3���D$�L$~8�S ����|#;D$}�L$ k�hFt��RxQP���҄�u�D$��;�|̊D$_^][��� ����������̃�SU�l$V�uW���Oh�   3�9\$(�D$�L$�t$�D$t�M0�L$$�6����t�\$��M0�L$$��q��;�~c�U�4���|I;t$}C�Gdi��   �L$(��RlQ�P���҄�u
�D$    ��|$ t�Gd���   Q�L$(��t����;\$|��|$ t�L$$�.6����t_^]�[��� _^]2�[��� ��j�hX�d�    P��(V�  3�P�D$0d�    ���   ����   �5�T$@����D��   �\$H����D{y�F<��|r;A}m�I�<� td���Rh�\$P�D$P���ҍD$P���D$<    诸����L$�\$(Q�L$D�[+���L$�D$8�����p��3��L$0d�    Y^��4� ��3��L$0d�    Y^��4� ��������������U����j�h��d�    P��(  SVW�  3�P��$8  d�    �]�CH�U;BD�F  �CX;BX�:  ���2  ;Ax�)  k�hAt�p���D$4u �K8;J8u����   ���Ѕ���  3��-3Ʌ�~'�x�d$ �C89�u�A����E��;P8t��;�|��T$4;J��  ��Ph�L$lQ���ҋu��Ph�L$|Q��Ǆ$D      ��j�L$pƄ$D  � ��� j �\$8��$�   �r ��� �L$<�\$,�'���L$T�'���D$4j j �D$DP�����$耩���D$,j j �L$\Q�����$�f�����T$T�T$LR�\$h�D$@P��$�   �vn����$���L$�$Q��Ƅ$L  膫����$�   Ƅ$@  �n���D$T���D$<��������Dz�T$�D$\���D$D��������Dz�T$�{T�G���w�$���3��
�   �����VT�J����d  �$����� ��t!����t���\$�d  ���\$�\$�U  ����u;�t���\$�?  ����t��u	�\$�*  ��$�   ��R���Ƶ��P�L$@�=���\$,��$�   P���)���P�L$X�=���\$,����Az�D$<�\$��   �D$T�\$��   �� ��   ����t�����\$�   ����u;�t���\$�   ����t��u	�\$�   ��$�   ��Q���!���P�L$@�=���\$,��$�   R��脵��P�L$X��<���\$,����Az
�D$D�\$�8�D$\�\$�.�����\$�\$� �� ����t����u�\$�
���\$��؍D$<P�L$Qj j�JK������t:�L$����   ���ĉ�L$0�H�L$4�H�L$8�H�L$<�H�L$@�H���ҍD$TP�L$Qj j��J������t:�L$����   ���ĉ�L$0�H�L$4�H�L$8�H�L$<�H�L$@�H���ҍL$|Ƅ$@   �l���L$lǄ$@  ������k�����$8  d�    Y_^[��]� 2���$8  d�    Y_^[��]� ���������������������������U����j�h��d�    P��h  SVW�  3�P��$x  d�    �L$ �E3�;ǉ��   ��  ;��   ��  i��   ��   �ȉD$0脸����;��t$$��  �D$\P�L$XQW��贻������  �T$LR�D$HPj��虻�����q  h��jj��$�   Q�s���D$DWW�T$|R���\$���D$p�$�������3  �D$DWW��$�   P���\$���D$x�$�������  �D$LWW��$�   Q���\$���D$p�$�e�������  �D$LWW��$�   R���\$���D$x�$�:�������  �M�|$4�|$8�|$<�|$@3�9<�t��   ����|�u�E��+�+ƿ   �D$�d$ ������   ����  �L$ ;AX��  k�h�ыJT�D@�3�ɋ+��ҋ@�X  ���P  �L$�1���u	�L$�1�;���   �ׁ�  �yJ���B�M������u��;���   ���W������^����t$ �U3���I �����t����   ;FH��   ����|ߋ|$$3�����   V���҉���   ����|�3�����   V���҉D�d����|�u�}3ۃ|�d ��   3������������   �T�;���   ���   +L����   hx�h\�h  h@��#����3���$x  d�    Y_^[��]� hx�h\�h  ��h��h\�h  �h̘h\�h  �h��h\�h+  땋T����u;�t�L��   +��T��#���u;�t;���   �   +L�9���   ����������E�]+ǉD$,��$�   +��|$(��3�+��Ӊ|$l��ɍt%�|$(ǋ|$,�<8���   �8 ��   �ɋ|$lu�΁�  �yI���A�|�d tD�F%  �yH���@�
��}�<� |)���u����hh�h\�hJ  �����<��u���������h����|$ �G(��9G,�O }P����3��hh�h\�hX  �Z�����$    �|$ �U������L$$�D4 tk�hGT�H@;HD�T4��   ����    t
�D4��   ��|3������|�d t�L4�L4�   ��wC�$���D$D���$j � �D$\��D$L���$j ��D$T���$j����   �ЉD�4�|�4���  �L$$���%  �yH���@���   P�҅�t�D4�����   ���҅����D4��	�M�<� u��|�U�<� u����   ���҃���������t$ �~L}�~L�N@}j�)���L$���9;ui�C��|��u\�C��|�|$ uN��L$t�T$x�� ���\$���$�   �P��$�   �H��$�   �P��$�   �H�ΉP�A���@(�L$�9{��   ��t��S�vh8�h\�h�  �s����C��|��uT�$�   ��$�   �� ���\$���$�   �P��$�   �H��$�   �P��$�   �H�ΉP�A���@(�L$�C9{ur��t�K�K�f�C��|�|$ t�C�S�$�   ��$�   �� ���\$���$�   �H��$�   �P��$�   �H��$�   �P�H���@���P(�S9{up�|$ t�C�C�a�|$ t��K�S�$�   ��$�   �� ���\$���$�   �H��$�   �P��$�   �H��$�   �P�H���(@���P(�S�   9F\}9F\�NP}P�Z+��3����    �|�4 ��   �E�<� t�~��  �yO���G����N��  ���yI���A�T$ �5�BD�U���ɍȋ������$�L$(�<ЋD�<j P�N����L$,PSW�@������XX�@8�M��u9t$ht5����P�E�   +�H���u�|$d t���P�P�E��+H�H�����)����t$ �Fh��9Fl�N`}P�+���F��9F�N}P�}����T$0Rj���A���D$T�X0�D$�D$D��$�   �X8�   ���P@�D$\�XH�D$L�XP�XX���������y�����\$��$�   �D$\�\$�D$l�$�%������\$�D$\��$  �\$�D$t�$��$������\$�D$d��$,  �\$�D$t�$��$������\$�D$d��$D  �\$�D$l�$�$���u��$�   �D$$�E+ƉD$p�D$4+ƉD$,�E3�+��D$4   �D$8   �D$<   �D$@   �D$0j,�Y������D$(��Ǆ$�      tjjj j��贁�����3��L$$Qj ��Ǆ$�  ������F���C�D$(%  �yH���@�@����   Pj���F�����  ��O��W���ZyK���C��Pl��t�D$L���\$�D$T��D$\���\$�D$d�$��W�|$$���H����L$l�<1 Pt%�T$0�2�L$ P����GDQ��Q���o���   �\$4�3�T$ k�h�D$tOTR�0RQ���m���L$,�1�L$(��  ��PTyI���A�|�d t	�@P   �A�@P   �3k�hWT�zP��~)3Ʌ�~#�zL�<��\$ i��   �[d���DP   ;JP|���j�P`j��Ph��ݐ�   ݘ�   �{R���\$(�D$$�����F����T$�B�L$ k�hAt��$x  d�    Y_^[��]� ������������������QUV�񍎐   �@_���L$3�;͉��   �l$u^3�]Y� �V8SW3�;�~�F4��    ;t
����;�|�;�|Q��趼����3�;�����W���C>���L$$�X�T$ �D$QRPS���9�����tiۨ   ��   _�\$��[^]Y� ��t�N4�W��    9V8u��|;~<�~8��i��   ��   j P��葧���K9��   u��|;��   ���   �D$_[^]Y� ��������V��F(W�|$P���-�������t7�NQ�����������t%�V,R���i�������t�F@�����$蒥����_^� ����������V��W�|$�F(P���͒������t2�NQ��蛓������t �V,R���9�������t��@V���'�����_^� ���������������j�h�d�    P�� SVW�  3�P�D$0d�    ���G8�\$@P���I�������t�O<Q���7��������X������؅�t|P����������tm�T$R���Y��P���D$<    �8����L$���D$8������\����t9�G@Pj���â������t%�OHQ���!�������t�GX�����$�J���������k����|6��t2��Rh�D$ P����P���D$<   �����L$ ���D$8�����U\���ƋL$0d�    Y_^[��,� ��������������j�h@�d�    P��$UVW�  3�P�D$4d�    ��L$�D$    ����|$D�E8P���D$@    ��������tl�M<Q���ސ������tZ�T$R���ː������tG�D$P���Ȓ������t4�M@Qj��蔐������t �UHR���"�������t�EXP���������L$�T$�D$�L$$�L$ �T$(�D$,�L$0���D$<�j����|E������=d��|7��t3�T$$R���>�������u �D$�L$�T$�D$$�D$ �L$(�T$,�D$0�L$�T$���ĉ�L$,�P�T$0�Hj �͉P�r���|$ t���g���L$$�T$(���ĉ�L$<�P�T$@�H�͉P��Y���L$$�D$< �Z���L$�D$<�����zZ���ƋL$4d�    Y_^]��0� ���U����j�hs�d�    P��   �  3ĉD$pSVW�  3�P��$�   d�    ��}���T$���T$�L$T�$�%���C8P���
���������   �K<Q�����������to�T$TR���qV��P��Ǆ$�       �����L$T��Ǆ$�   �����Y����t5�C@P��訟������t#�KDQj��脟������t�SLR��聟�������CPtP���o��������CTt1P���]�������t"�CXP���K�������t�K`Qj���G��������mh����}0����   �T$<R�������������   �D$<P���ݠ���   ��t8��Rh�D$,P����P��Ǆ$�      �����L$,��Ǆ$�   �����X��3��ˉD$h�D$l�D$p�D$t�D$x�D$|�+T���������D$ht�L$hQj���@��������D$h tG�T$hRj���&�������t4݃�   �����$��������t݃�   �����$�ҟ������Ƌ�$�   d�    Y_^[�L$p3���  ��]� ��������V��FW�|$P����������t�NQ���;��������N$tQ���ɝ������t�V(R��距����_^� ���������������V��W�|$�FP��荌������t�NQ��������3Ʌ��L$t�T$R���b����L$����w)�$�<��F$    ��F$   ��F$   ��F$   ��t��(V��������_^� ���
�������V��FW�|$P��������t9�NQ���>�����t*�V,R���Ϝ����t�F0P��远����t�N4Q��谜��_��^� ��������V��W�|$�FP��荋����tW�NQ��������tH�V,R���o�����t9�F0�L$Q�ωD$�W�����t!�|$ ���V0��4V�=����> }�    _��^� ����������j�h��d�    P��   �  3ĉD$|SUVW�  3�P��$�   d�    ��$�   ���t$H�   ��    ���������y�G8P��越��������   �O<Q��蠊��������   �L$(����T$(R��Ǆ$�       腌������tN�L$(�T$,���ĉ�L$@�P�T$D�H�ωP��P���L$(�T$,���ĉ�L$@�P�T$D�H�ωP�PT���L$(Ǆ$�   ������T����tL�G@P�����������t:�ODQj���ى������t&�WL�D$P�͉T$�Ή������t�|$ ���OL3����D$�Xt�T$R��裉�����D$;�w.�$���GP    ��GP   ��GP   ��GP   ��_P3����D$t�D$P���T������D$��w@�$� ��GT    �0�GT   �'�GT   ��GT   ��_T��GT   ��GT   ��t"�OXQ�����������t�W`Rj������������c�����  ������=d���  �D$P���DP����Ǆ$�      tC�L$Q��詊������u0�T$8R���P����L$�P�T$�H�L$ �P�L$8�T$$�RS��3�2ۅ��D$x�D$|��$�   ��$�   ��$�   ��$�   t:�D$xPj����������t%�|$xu��L$xQj����������t���_���T$�L$���ĉ�T$0�H�L$4�P�H���R���L$Ǆ$�   �����R���&��tN�T$HR��菈������t=�D$`P���|�������t(���   Q����������t�Ǹ   W����������Ƌ�$�   d�    Y_^][�L$|3����  �Č   � ��ȲѲڲ���!�*�3�8�A�����QS�\$W��j h � @�ˉ|$�9������tnVj j��袝��������|$tW���̗����U3��t*3�;l$}"��t�D$�H�9�B �S�Ћ�����H��u؋�������]u	^_3�[Y� ��^_[Y� ����������QS�\$W��j h � @�ˉ|$�u8������tqVj j������������|$tW���,�����U3��t-3�;l$}%��t�D$�H�9�B �S�Ћ������   ��uՋ��������]u	^_3�[Y� ��^_[Y� �������QS�\$W��j h � @�ˉ|$��7������tnVj j���b���������|$tW��茖����U3��t*3�;l$}"��t�D$�H�9�B �S�Ћ�����h��u؋��A�����]u	^_3�[Y� ��^_[Y� ����������QS�\$W��j h � @�ˉ|$�57��������   Vjj��辛��������|$tW��������U3��t-3�;l$}%��t�D$�H�9�B �S�Ћ����Ǩ   ��u�3��t+3�;l$}#�L$�Q�D:8P��耗�������Ǩ   ��u׋��i�����]u	^_3�[Y� ��^_[Y� �̃�SUVW�|$j��j��������3�;��  W�M�b�����;��  W�M �N�����;���  W�M0�ʻ����;���  W�M@�������;���  W�MP������;���  W�M`�a�����;���  W�Mp�������;���  W���   �x�����;��  ���   P���p�����;��f  ���   Q���W�����;��M  ���   Sh � @�ωT$�u5����;��+  �\$�\$���D$9D$}T���X����t���   �T$���   �3ۅ�����P�ّ������t��tS���_�����D$�D$�   ��u����˾������   3�;���   Sh � @����4����;���   �\$�\$���$    �L$9L$}T���?X����t���   �D$���   �3ۅ���Q���9�������t��tS���_�����D$�D$�   ��u����+�����t��t���   R���%�����u3�_��^][��� ��̃�8�D$<SU�hh��@xVW�l$�D$~U3ې�D$L�pd󍾀   �������u)��诚����t�L$Q��������   �L$�L�����   ��u��D$��~h3�D$�d$ �T$L�rt��^0���-����u=3�9~~6���F����|";D$}�L$Li��   �Qd���   P���O����;~|̃�h�l$u�_^][��8�����������j�h?�d�    P��   SUVW�  3�P��$�   d�    ���|$3���$�   �t$ �t$D�t$d�t$,�t$|�K����$�   �D$ P�͉�$�   豀���؄�t2�L$DQ��蟀���؄�t �T$dR��荀���؄�t�D$,P���{����ظ   9D$ |9D$D|9D$d|9D$,}2��:��t6�L$|Q���H����؄�t$���   R�������؄�t�Ǩ   W��� ����؋|$�D$,��9G}P���w���ۉt$��   �D$,9D$��   j(��������D$X��Ƅ$�   t���������3���B$U��Ƅ$�    �Ѕ������W����u&j ��������L$(Q�ωD$,蹘����Bj������L$(Q�ωt$,蜘���D$���e����|$�W�D$D�� 9G�T$p}P���@v�����D$    ��   �D$D9D$��   j(�+������D$X��Ƅ$�   t����������3���B$U��Ƅ$�    �Ѕ����������u&j �������L$(Q�ωD$,������Bj������L$(Q�ωt$,�җ���D$���e����|$�w(9w\�OP�t$(}V�L��3����D$~��tP���&&���D$��;ƉD$|�D$ ��09G}P���Cu�����D$    ta�T$ 9T$}Wj@�6������D$X��Ƅ$�   t���\�����3���P$U��Ƅ$�    �҅��D$0P���Ét$4�����D$��u��t$,3�;��D$4�$�|$8�|$<�|$@~F}�t$<VW�L$<��$;ǉD$8t$�L$@;�~��+���R��WP���  ���t$@��|$@�|$<�t$,;�Ƅ$�   �D$H�$�|$L�|$P�|$T~F}�t$PVW�L$P��$;ǉD$Lt$�L$T;�~��+���R��WP�i�  ���t$T��|$T�|$P�L$�D$ ���   9AƄ$�   }P�W���L$�D$d��p9A}P����L$�D$,��`9A}P����ۉ|$h�~  ��;D$ �  �L$3�P��$�   �t$`��&���ۋ���$�   t �L$Q���s|���؄�t�T$R���a|���؄��G0�D$tta�L$tQ���G|���؄�tO9t$t��$�   ��P�͈W0�(|���؄�t0�OHQ����|���؄�t��`W����|���؄�t�T$\R����{���؃|$\}2ۄۉt$`��  �D$\9D$`��  3��ۉ�$�   tD�L$Q���{���؄�t��$�   R���{���؋�$�   ���t;�t��������������   ��   ��t*��$�   Pj���m{���؄�t��$�   Qj���V{���؄ۉ|$lt�T$lR���0{���|$l��}2ۋ�$�   �L$PV�$���ۉD$X�|$$��  �I �L$$;L$l��  �L$�Ah�T$XPRj �>T�����~8W�L$8�Op����t�D$P���z���؋;L$th��h��hM  ht��L�������t�T$xR���z���؍D$xP�L$L��o�����D$ t;�L$Q���x���؄�t�V@R���Sz���؀|$ t�F@����   ;D$(��   �����   ;D$p��   �ۉF<�FL�D$0tk�L$0Q���z���؄�tY�|$0 ��$�   ��P�͈VL��y���؄�t9��$�   Q����y���؄�t$���   R���Mz���؄�t�ư   V���9z���؃D$$��������GhD�h��hZ  ht��F@�����(���� h�h��hb  ht������F<������2ۃD$`���g����D$h���ۉD$h������L$�(�����  3�3��D$���    ;D$ ��  �L$i��   ��   �T$R�͋��(w���|$ t>�D$$P�͉|$(��Z���L$$��Q���a�����;ǉ��   u�L$$;�t	��Bj�ЋD$���ۉD$u��"  ���V����|$3�9t$,�t$�   �I �D$8����|;Oh|_�T$L�����D$x|;Gh|K�Wdi��   i��   �Q@��|;T$p�|$}�x@ }�P@��@@��|;D$p�|$}��}�A@�t$��;t$,�t$|�3�9Gh�D$~U���$    �Oi��   Gd���F<��P���D`���F@��|;D$(}�WTk�h��8V�LH�$m���D$��;Gh�D$|����"��j ���4�����R�����z���I�����uQ3�9|$ �D$~=��L$��i��   ��   ���   ;�t��Bj�Љ��   �D$��;D$ �D$|Ą���   ��$�   ��   3��ۉD$�   3�;D$ }s�L$i��   ��   �T$R�͋��u���|$ t=�D$$P�͉|$(��X���L$$��Q���T�����;ǉ��   u�L$$;�t	��Bj�ЋD$���ۉD$u����uJ3�3�9|$ �D$~<�l$��i��   ��   ���   ;�t��Bj�Љ��   �D$��;D$ �D$|ȋ|$W��������u$h̙h��h�  ht����������|$�   9t$|u���������t���   3�9t$T��$Ƅ$�   �|$Ht �D$L;�tVP�L$P��$�t$L�t$T�t$P9t$@Ƅ$�    �|$4t �D$8;�tVP�L$<��$�t$8�t$@�t$<��$�   Ǆ$�   �����T@���Ë�$�   d�    Y_^][�ļ   � ������V��F�V;�uS����Ɂ�   v��|��q ;�}�������   ��;�}BP�������N�F�Ƀ��N��^Í��F�Ћ�Bj �ЋF�V����P���z����N�F�Ƀ��N��^�������V��F�V;�uN��k�h��   v��|�C� ;�}�������   ��;�}=P���	���N��k�hF���N^�k�hFj ��ȋB�ЋNk�hNQ��������N��k�hF���N^�V��F�V;�u@��iɨ   ��   v��|��0 ;�}�������   ��;�}2P���5
���(i��   Fj ��ȋB�ЋNiɨ   NQ�������N��i��   F���N^�����̃�UVW������l$(3��D$P�L$Q�͉t$�t$$�t$(�t$�t$�t$ 脻������   �|$ � @Suf�T$R�D$P��� ����؄�tQ�|$uH�L$Q���s���T$R�ϊ�����9t$~*�I ��t#��������ȋB$U�Ѕ��Ã�;t$|��2ۋ��B�����u[_^��]��� ��[_^]��� _^��]��� �������̃�UVW�������l$(3��D$P�L$Q�͉t$�t$$�t$(�t$�t$�t$ 蔺������   �|$ � @Suf�T$R�D$P�������؄�tQ�|$uH�L$Q���r���T$R�ϊ�����9t$~*�I ��t#���u����ȋB$U�Ѕ��Ã�;t$|��2ۋ��R�����u[_^��]��� ��[_^]��� _^��]��� �������̃�UVW�������l$(3��D$P�L$Q�͉t$�t$$�t$(�t$�t$�t$ 褹������   �|$ � @S��   �T$R�D$P�������؄���   �|$��   �L$Q���q���T$R�ϊ����9t$�t$,~h�I ��ta���C������P$U���҅��Ä�t0�G��9F8t%h�hؚh�  ht��l����O�����N8�D$,��;D$�D$,|��2ۋ�������u[_^��]��� ��[_^]��� _^��]��� ���������̃�UVW���S���l$(3��D$P�L$Q�͉t$�t$$�t$(�t$�t$�t$ �d�������   �|$ � @Suf�T$R�D$P��������؄�tQ�|$uH�L$Q����o���T$R�ϊ����9t$~*�I ��t#���%�����ȋB$U�Ѕ��Ã�;t$|��2ۋ��"�����u[_^��]��� ��[_^]��� _^��]��� �������̃�UVW������l$(3��D$P�L$Q�͉|$�|$$�|$(�|$�|$�|$ �t�������   �|$ � @S��   �T$R�D$P�������؄���   �|$��   �L$Q����n���T$R�Ί��M���D$��~*��I ��t!��������ȋB$U�Ѕ��D$�Ã�;�|ۃ|$|83�;�~2�|$,��t*�N�T$,�D8P���p���D$,�   ��;|$��|��2ۋ�������u[_^��]��� ��[_^]��� _^��]��� �����������j�h��d�    P��DSUVW�  3�P�D$Xd�    ��\$h�D$$P�L$,3�Q�ˉl$0�l$,�Ȅ����;��~  �D$(��u�T$$RS���������`  ���W  S�N�}�����;��F�D$tS�N �f�����;��N(�L$,tS�N0������;��V8�T$��  S�N@�������;���  S�NP�������;���  �FX����   �l$ �~T|$ �G<���w`��   ;D$,��   ���3���؍D$HP���4����Rh�D$8P���D$d    �ҋL$H�T$L���ĉ�L$`�P�T$d�H�N$�P�G<��R���D$t��N����t���nD���L$8�T$<���ĉ�L$P�P�T$T�H�ωP�6���L$8�D$` �i7���L$H�D$`�����X7���\$h�D$ h��;nX����S�N`����������  3�9nh�l$ ��   �~d�D/<������   ��   ;D$��   ���2���؍D$8P���3����Rh�D$HP���D$d   �ҋL$8�T$<���ĉ�L$P�P�T$T�H�N�P�G<��R���D$t��M����t���dC���L$H�T$L���ĉ�L$`�P�T$d�H�ωP�5���L$H�D$`�_6���L$8�D$`�����N6���\$h�D$ �����   ;Fh�D$ ����S�Np�����������   3�9Fx~3ɍd$ �Vt�t`����h;Fx|�S���   ��������ts3�9��   ~;3����   �D9,υ����   |;D$}�V4��P�XO�����Ǩ   ;��   |Ǎ��   Q�L$l�k������t�L$h���   R�pk�����\$h3�V�q�����;��  �|$$��  ���   �L$0Q�T$$R�ˉD$4�l$(�l$8�l$<脲����;���  �|$  � @t3��   �l$3ۋD$;D$,��   �l$h�L$Q���Dh������t]�|$ tV�T$R���D$     �L�����D$��t8���   P��j������   ���   �����    u�L$��t	��Bj�ЃD$�è   ���k����\$h3��� �����u3��  ;��  �L$0Q�T$$R�ˉl$(�l$8�l$<萱����;���   �|$  � @t3��   �l$3ۋD$;D$,}{�l$h�L$Q���Tg������tQ�|$ tJ�T$R���K�����   ���D$P�膫�����   ���   �����    u�L$��t	��Bj�ЃD$�è   ���{����\$h3��������u3��5;�t1�|$$|*�L$h���   S�yh�������|��|�    �\$h3������=
1��}���   �L$Xd�    Y_^][��P� ��̸������������̋L$h��2����   � ���������̸������������̋D$V��;�t,�H�N�P�V�H�N�P�V�H�N�PP�ΉV�S����^� ���V�t$Wj j��h � @�������u_3�^� �GSP���x���؄�t/�OQ���px���؄�t�WR���_x���؄�t�GP���Nx���؋��5�����u2���[_^� �����̃�V�t$3�W�D$�D$���D$P�L$Qh � @���u�����u
_3�^��� �|$S�Ä�t@�WR����f���؄�t/�GP����f���؄�t�OQ���f���؄�t��W���f���؋��#�����u2���[_^��� ̸p������������SU�l$��;�t@�E�C�M�C�@�K�UV�K�SW�UR�ЋM$�K$�u(�{(�   �U���R��_^]��[� �������������V�t$Wj j��h � @�������u_3�^� �GSP����v���؄�t/�O$Q����v���؄�t�WR���/{���؄�t��(W�������؋�襡����u2���[_^� �����̃�V�t$3�W�D$�D$���D$P�L$Qh � @��������u
_3�^��� �|$S�Ä�t@�WR���Oe���؄�t/�G$P���>e���؄�t�OQ���l���؄�t��(W���f���؋�蓣����u2���[_^��� ̋Q2���t%�I��~V�t$��t��~Vj(QR�h*�����^� ��������������̋Q2���t%�I��~V�t$��t��~Vj(QR�*�����^� ��������������̋D$�L$�����PQ�������� ��j�h��d�    PQV�  3�P�D$d�    �t$�t$���D$    t/����B������F�F�F3��@��F    �F     �F�F�L$d�    Y^��� ��������j�h��d�    P��HSUVW�  3�P�D$\d�    �����   ���   �l$ �D$�~��P�7�������D$(��   �틈�   �L$$��   �D$    �l$���   t$�^(���W.��3�9n~l�V����|Z;D$}T���   ���D���|C;D$$}=�T$(i��   ��   �L$,Q���=���P���D$h    �=1���L$,�D$d������-����;n|��D$`�l$�i����l$ �|$ �\$l~ �l$3����   S��aB����(��u�l$ ��~3����   S��AB����`��u�   �L$\d�    Y_^][��T� ��������������j�h�d�    PQV�  3�P�D$d�    j(�Gv�������t$���D$    tB���@������F�F�F3��@��F    �F     �F�F�ƋL$d�    Y^���3��L$d�    Y^����������������j�h;�d�    PQSVW�  3�P�D$d�    ��j(�u�������t$������D$    t.���@��3��@��^�^�^�F    �F     �F�F�3����\$t0;�t,�G�F�O�N�W�V�G�F�O�N�WW�ΉV��L���ƋL$d�    Y_^[�����������������VW�|$��t5h������A����t%�t$��th������A����tW�������_�^�_2�^�������������V���@��G���D$t	V�v������^� ������������VW�|$��t5hp����ZA����t%�t$��thp����BA����tW������_�^�_2�^�������������QU�l$Vj ��jh � @�͉t$�����t]�FSWP�͉D$��p����3���t-3��d$ ;|$}!�D$�H�1�B �U�Ѕ��Ã���(��uً�袛����u_[^]Y� _��[^]Y� ������������SVW���G�4���3��9_~&U3���I �G�(�(�B�Ѓ���(;_�t�|�]_��^[�������������QU�l$Vj ��jh � @�͉t$�����t]�FSWP�͉D$�p����3���t-3��d$ ;|$}!�D$�H�1�B �U�Ѕ��Ã���`��uً������u_[^]Y� _��[^]Y� ������������SVW���G�4@3���9_~)U3����    �G�(�(�B�Ѓ���`;_�t�|�]_��^[�������������V�t$Wj j��h � @��������u_^� SV�������؄�tV�O������؋�������u2ۊ�[_^� ��VW����>���NX��~3��VT�t`��h��u�Nh��~3��I �Vd���   �   ��u�Nx��~3��I �Vt�t`��h��u񋎈   ��~3���I ���   ���   �   ��u�D$P�����;��P���b<������t[h�����`>����tK���   ��tA�P�҉p ~3ɍ�    �p�D ��(��u�P��~3����    �p�D1X��`��u�_^��������������SV��^��xUW�<�����N�9�P�j �ҋF�3ɉ�H�H�H�H�H�H�H�H �H$�F�P���J�������(��}�_�F    ^[������S�\$��UVW��}N3�9nt:�~��x!����ۋN��P�U�҃���(;�}�N��PUQ���҉n_�n�n^][� �F;�}x�N��PSQ����3�;ǉFtT�V��+ʍ����Q����WP�G�  �F��;�}"�<������+�N�Q���s�����(��u�_�^^][� �~�~_^][� ~V���;�|'�<���+������N�9�B�j �Ѓ�(��u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� �����U�l$V��;��~   �ES3�;��^[��^]� 9F}P����9^t�E;ÉF~�W3��E�N��;�t*�P�Q�P�Q�P�Q�P�Q�P�Q�PP�Q�F������(;^|�_[��^]� ��^]� �����������SVW�����   �K������ˋ���������k	��_�^[�����̋D$P���   ������� ����������j�hs�d�    PQVW�  3�P�D$d�    ��t$��8��3�����|$�F�$�~�~�~ �N(�D$�Y$������F�F$3��~X�F�F�ƋL$d�    Y_^����j�h��d�    PQSVW�  3�P�D$d�    ���|$����O(�D$   �$��3�9_ �w�\$��$t�F;�tSP����$�^�^�^���D$������?���L$d�    Y_^[���UW��3�9o�x�t>V�w��x#S����ۋO��P�U�҃���(;�}�[�O��PUQ���҉o^�o�o_]��������̋D$��S�U�V�t$�PV���c���������t)��t%;�t!W3�9{~����B���Ѓ���(;{|��_^][� �����������V��V2���tQ�N��~JW�|$��t@��~9Wj(QR����3���9~~%S3����    �F���B�Ѓ���(;~|�[�_^� ���������������V��V2���tQ�N��~JW�|$��t@��~9Wj(QR�u��3���9~~%S3����    �F���B�Ѓ���(;~|�[�_^� ���������������V��F�V;�uS����Ɂ�   v��|�;33 ;�}�������   ��;�}BP��������N�F�����N��^Í��F�Ћ�Bj �ЋF�V����P��������N�F�����N��^�������V�������D$t	V�m������^� ��j�h��d�    PQ�  3�P�D$d�    �L$�L$���D$    t�V����L$d�    Y��� ����j�h��d�    PQ�  3�P�D$d�    j`�j�����D$���D$    t��������L$d�    Y���3��L$d�    Y���������������j�h+�d�    PQVW�  3�P�D$d�    ��j`�j�����D$���D$    t���������3����D$����tW���P����ƋL$d�    Y_^���������������V��������D$t	V�k������^� ���؛�5�������̃�UVW���s����l$�D$P�L$Q3�h � @�͉t$�t$�t$ 軟����th�|$S�Ä�tC�T$R���.U���؋D$P������9t$~#��t���_�����ȋB$U�Ѕ��Ã�;t$|݋��p�����u
[_^]��� ��[_^]��� ������j�ha�d�    P��SVW�  3�P�D$d�    ���_��xU�4[���O�1�P�j �ҋGj`�j P�̨  �O��ΉL$�L$�D$     t���������`���D$ ����}��G    �L$d�    Y_^[����S�\$��UVW��}K3�9nt7�~��x����N��P�U�҃���`;�}�N��PUQ���҉n_�n�n^][� �F;�}{�N��PSQ����3�;ǉFtW�V��+ʍI�R��Q���WR��  �F��;�}&�<@����+荤$    �F�P��������`��u�_�^^][� �~�~_^][� ~S���;�|$�<@+�������N�9�B�j �Ѓ�`��u�9^~�^��F�RSP�Ή^��3�;��Fu�N�N_^][� ��������U�l$V��;�tX�ES3�;��^[��^]� 9F}P����9^t�E;ÉF~�W3����E�N�P�� �������`;^|�_[��^]� ��^]� �����V���؛�"����D$t	V�uh������^� ������������UW��3�9o���t;V�w��x S�v���O��P�U�҃���`;�}�[�O��PUQ���҉o^�o�o_]�����������̋D$SU�@V�t$��PV���f���������t)��t%;�t!W3�9{~����B���Ѓ���`;{|��_^][� ��������������V��V2���tQ�N��~JW�|$��t@��~9Wj`QR����3���9~~%S3����    �F���B�Ѓ���`;~|�[�_^� ���������������V��V2���tQ�N��~JW�|$��t@��~9Wj`QR�u��3���9~~%S3����    �F���B�Ѓ���`;~|�[�_^� ���������������V��F�V�@��;�uJ��   v��|�]U ;�}�������   ��;�}<P���7����N�I��F���N^�Nj ��B�ЋF�@��NQ���C����N�I��F���N^����������������V�������D$t	V�f������^� ��V��� ������D$t	V��e������^� �����������̃�UVW��������l$�D$P�L$Q3�h � @�͉t$�t$�t$ �������th�|$S�Ä�tC�T$R���nO���؋D$P���0���9t$~#��t��������ȋB$U�Ѕ��Ã�;t$|݋�谍����u
[_^]��� ��[_^]��� ������j�h��d�    PQV�  3�P�D$d�    ��t$�N�D$    � ��������D$�����؛�m����L$d�    Y^���������������VW�|$��;�tVW�>����G�N;�tP����3�9F~3���I �V�t
 ����(;F|�3�9F~3���I �V�t
X����`;F|�_��^� ������̃�VW�|$��D$P�L$Qh � @���D$    �D$    �o�����u_^��� �|$S�Ä�tXW���^�����3�9F~3ɍI �V�t ����(;F|��t,W�N�������3�9F~3ɍ�    �V�t
X����`;F|��������u2ۊ�[_^��� ������j�h��d�    P��V�  3�P�D$d�    ��t$�Q���3��,����   ���   ���   ǆ�   ��D$$���   ���   ���   ǆ�   ��   �D$$�F(�D$P����B+����N�P�V�H�N�P�V��/�F��/�N��/�V ��/�F$�ƋL$d�    Y^�� �������j�h��d�    PQV�  3�P�D$d�    ��t$�,����   �D$    �?������D$���������L$d�    Y^������������������V�������P� �����   �D$��P���   �������^� ��j�h+�d�    PQ�  3�P�D$d�    h�   ��_�����D$���D$    t���;����L$d�    Y���3��L$d�    Y������������j�h[�d�    PQVW�  3�P�D$d�    ��h�   �a_�����D$���D$    t����������3����D$����t;�tW�������Ǹ   W���   �g����ƋL$d�    Y_^������VW�|$��tKh������+����t;�t$��t3h������+����t#;�tW�������Ǹ   W���   � ���_�^�_2�^�������V��������D$t	V�`������^� �̋D$= �  r= �  r=�� v3�ø   ��������������̋L$��w�D$��   Á��  w�D$���������?�ɀ��H�   Á���  w+�D$��������������?�ʀ��?�ɀ�P�H�   Á��� w9�D$��������������?�ʀ�P������?�ʀ��?�ɀ�P�H�   Á����wV�  ���+�������ЋD$����������?�ʀ�P������?�ʀ�P������?�ʀ��?�ɀ�P�H�   Á����wU�D$��������������?�ʀ�P������?�ʀ�P������?�ʀ�P������?�ʀ��?�ɀ�P�H�   �3������U�l$V�����x���E ^�   ]ÊЀ�����u8���;  �I�р��������'  ��?��ȃ�w�^�M �   ]ÊЀ�����uR����  �Q������$�<���  �I��?����$��<���  ��?��ʁ��  w�^�M �   ]ÊЀ�����uo����  �Q������$�<���  �A��?��֋�Ѐ������n  �I��?���р��ƀ���U  ��?��ȁ���  w�^�M �   ]ÊЀ�������   ���   �Q������$�<��  �A��?��֋�Ѐ�������   ��?��Ƌ��A�Ѐ�������   �I��?���р��ƀ����   ��?��ȁ��� w�^�M �   ]ÊЀ�������   ����   �Q������$�<�ux�A��?��֋�Ѐ�����ua��?��Ƌ��A�Ѐ�����uJ��?��Ƌ��A�Ѐ�����u3�I��?���р��ƀ��u��?��ȁ����w�^�M �   ]Ã^3�]��������������̋D$= �  s�L$f��   �= �  rF=��  w�T$f��   �=�� w+�L$-   ����
%�  �� (  - $  f�Af��   �3����������UV�t$��W��   �|$����   �l$����   �f�� ���   f�� ���   ��|4f�� �s-�Ff= �r#f= �s�Ɂ���  ����
_�^�M �   ]ËD$����   �H�����Su]�XS���������tM�   ;�~<�I �Ff�� �r.f�� �s'�P;�}f�� �s�LFf�� �rf�� �r��;�|ǉ] [_^]�[_^3�]���_^�U �   ]ËD$��t�_^3�]���������Q�L$��SW�=  �|$���1  �\$���%  ��Q�D$�T$�D$ (  f=���   ��|If�D$f= �s>�Q�T$	�Q�T$�T$�� $  f���w�L$��-��  ��
��_�   [YËD$����   �P�����U��   �hU��������tq�   ��;�~^V��T$�Q�T$�T$�� (  f���w<�p;�},f�|$ �s#�Q�T$�Q�T$f�T$f�� �rf�� �r	�ƃ�;�|�^�+]_[Y�]_3�[Y��D$�_�   [YËD$��t�_3�[Y���̃�0�  3ĉD$,�T$H�ҋL$@�D$TS�\$<W�\$�L$�T$�D$(t�    �|$D���u����  3�f9;t
��f�<{ u�����  ����  �|$L u�D$    �D$L��������  3�9D$<t(��~$�f����u���f����u�   +����\$�L$TUV3��L$(�L$`3�;Ɖt$$�L$,ty����   �T$R�D$(P��+�Q�sR���������D$ ��   �L$�D$4PQ�����؋D$ ����t�+;T$T��   S�L$8Q�P��  ��t$ �;��\$|��~��~~���    �T$R�D$(P��+�Q�sR���������D$ ~O�L$�D$4PQ�����؋D$ ����t�+;T$T!S�L$8Q�P�
�  ��t$ �;��\$|��	�\$�L$$�T$�D$��t
;l$T}�( �D$0��t�s���t�D$$�^��]_[�L$,3����  ��0Å�t�
��t��L$4_[3�3��ڐ  ��0������������̋T$����t�    U�l$W�|$ ���u���^  3�f9} t��f�|}  u����C  ���;  �|$( u�D$$    �D$(�����|$$ �  3�9D$t%��~!�M f����u���f����u
�   +����L$0SV3��L$�L$<3�;Ɖt$�L$tH;���   �T$(R�D$P��+�Q�Tu R��������~i�L$,��t;\$0}V�T$(�����;�|��I;�~I�D$(P�L$Q��+�R�Du P�!�������~%�L$,��t;\$0}�T$(�����;�|���L$�T$4�D$,��t;\$0}��    �D$@��t�Lu ���t�D$�^��[_]��Å�t�
�D$8��t�(_3�]������������������̃�SU�l$��V�j  �t$ ���^  �\$(���R  �E ��x��^�]�   [��ÊȀ�����u9��|4�M�р���������   ��?��ȃ���   ^]��   [��ÊȀ�����uc��|^�M�р���������   ����?��E�Ѐ�������   ��?���=   ��   = �  v= �  r}^�]�   [��ÊȀ�����ue��|`�M�р�������uO����?��E�Ѐ�����u9����?��M�р�����u#����?ȍ�  ��=�� w^]��   [���W�L$Q�|$$�Ƌ��D$$    �D$���������L$$������~)��u%�T$�� �  r��  ��=� w_��^]�[��ËT$�\$(����  �{	��#�;���  ��m�{W�   ��������tN�t$$;�~@�d$ �)��y5�Ѐ�����t+�Ѐ�����t!�Ѐ�����t�Ѐ�����t$�<�t��;�|ċD$,�8_^]��[���R��������t��u�L$,_��^]�[��ËD$$;���   �� (�����  ��   ��t	����   ��   ��   �T$R+ƍ.�|$$�D$�����������������   �D$ ��t��uxf�D$f�L$j j j �T$,Rjf�D$,�D$$Pf�L$2j�L$4Qj �D$D    �D$4�����2�����$��u,�|$  u%�L$Q���������t�T$,�7_^�
�][��Ë[S��������t�D$,_���^][���_^]3�[���^]3�[�������������̋T$��VW3�;�t�:�t$$����D$ u;��
  3��8 t�I ���<0 u�;���   ;���   9|$,u�|$(�D$,����
9|$(��   �L$4S�L$�L$<3�;��|$�L$~{U�T$R�L$Q��+�R�P����������~Q�T$�L$,QR��������|$0 t%�;L$4*��f�T$,�L$0f�Yu
f�T$.f�TY؋D$(�;�|��	�L$�D$(�T$8]�L$,��t;\$0}f�Y  �L$@��t��9��t�D$���[_^���;�t�
�L$<;�t�_3�^�������������������������U����j�h��d�    P��h  SVW�  3�P��$x  d�    �}��$�   P���D$/ �A���]��$�   Q���A��j ���<A��P��$   Rj ���*A�����S���jj�L$\趮��j �L$XǄ$�      �Ч������$�   P��Q�������$�   R��P�|����\$D��j�L$X蚧���D$4j�X�L$X舧����$�   Q��$�   R���A��������j �L$X�_����j �X�L$X�O���j�L$X���B����@�����Aujj �L$\虧���D$,   ��D$,    j�L$X�����@��j��4�L$X�\$8�����@��$�   ��P��4��$�   Q�\$D������$  ݜ$�   R��$�   P��������ݜ$�   �D$<��$�   Q��$�   R���L$d�$�c������  S���D$/������t�E���t��E����  ���  �CP���������t�E��t����E����  ����  �wS���������t�E��t����E����  ����  �CP��������t�E���t��E���i  ��d  ��D$DP��$�   Qj���L$h�$�T������D$+�8  �E���L$,t�D�D��E��t��    �t$L+���݄$�   ���\$4����A��   �4�    �D4D����$�   �$P���?���L$L+������$�   �$R����>����$�   P��$�   ������T$,�D$4��������   ��;����A��   ��$�   Q��$  R���i@����$�   P��$0  Q���R@����$,  R��$�   �����\$<��$  P��$�   �v����D$<�(J���D$,��������Au9���D$+ ���؍L$TǄ$�  �����\����D$+��$x  d�    Y_^[��]���������Au��D$+ ������$P�\$�D$�HQ�L$�PR�T$P�D$$�@x������`�\$��`�A��`���\$�B���$PQR�|���������<���3�V���F�F�F�N �F�F�F�F�D���N$�D���N(�D���N,�D���N0�D���N4�D���N8�D���N<�D���N@�|D���ND�tD���NH^�kD�������������V�t$Wjj��h � @���������>  SW���H���؄��  �GP���F���؄��  �O Q���I���؄���   �W$R���I���؄���   �G(P���I���؄���   �O,Q���nI���؄���   �W0R���YI���؄���   �G4P���DI���؄���   �O8Q���/I���؄�ts�W<R���I���؄�tb�G@P���I���؄�tQ�ODQ����H���؄�t@�WHR����H���؄�t/�GP���*E���؄�t�OQ���E���؄�t�WR���E���؋���o����u[_^� ��[_^� ������������̃�SVW�������|$�D$P�L$Q3�h � @�ω\$�\$�~�����N  �|$�+  9\$�!  V���5���؄�t@�VR���y3���؄�t/�F P���X8���؄�t�N$Q���G8���؄�t�V(R���68���؃|$��   ����   �F,P���8���؄�ts�N0Q���8���؄�tb�V4R����7���؄�tQ�F8P����7���؄�t@�N<Q����7���؄�t/�V@R����7���؄�t�FDP���7���؄�t�NHQ���7���؃|$|7��t3�VR���2���؄�t"�FP���2���؄�t��V���u2�����2ۋ���p����u	_^[��� ��_^[��� j�h)�d�    PQV�  3�P�D$d�    ��t$�N �B���N$�D$    � B���N(�D$��A���N,�D$��A���N0�D$��A���N4�D$��A���N8�D$�A���N<�D$�A���N@�D$�A���ND�D$�A���NH�D$	�A�����D$
�����ƋL$d�    Y^���������������S�\$��Wt)�|$��v!VW�_��������tWSV覉  ����^_[�_3�[��������̋D$�� Wt;��t.��t"hԝhĝh�   h��賠����2�_� �9�A��y�A�3�3�S�\$��U�l$Vr|��sb���ދӃ� ��;�w+r;�s%h|�hĝh�   h���T�����^][2�_� �ËЋ�;qu;Qt�q�Q�A    ^][�_� ��|���vҋ�����;�w�r;�w�h(�hĝh�   h��������^][2�_� ���������������QSU�l$W�}���ى\$�B  V��    �w�;ƋW�  �K;��  ;U��   r	;u ��   �G;ЋOr'w;�r!h �h�h�  h���X������   � t
+�ً��3�3�S R�]����3���F�F�F�F�F����F�Fw��v�F �F�OSQP謇  ���\$�{ u�s�S��C��t�p�s�G�F�O�N�W�V�G�F�D$��@�v;�wr;�r�ʋƋl$��C���������h �h�h�  h���y�����^�E;C�Mwr;w�K�C_][Y� ������̃�����Q�$�T$u$��u 9Qt2���� �y u�y ����� �A��tރ8 u�U�i��t�} t	2�]��� VW3��D$    3�S��$    ;8uo��t�O;Huc�W;Pu[�H�x;ϋP�XrKw;�vE9\$u?;�u;+�ϋ|$��;�w+r;�s%���@���T$��u�;�u�t$;�wr�D$;�s[_^2�]��� �D$;ur�w;Ev�;uw�r;Ew�[_^�]��� ��������̃�SU��]3��ۉD$�D$��  VW��D$�S;S�K�\$r(w;Kv!h`�hL�h%  h���ݜ������   ��u��u��t;h�hL�h2  ��p;�u�@;�th��hL�h=  h��葜�����s+s�{{��u%��u!h��hL�hF  h���a������   ��L$��D$;Er<w;M v5;]u�{ thP�hL�hP  h���������u +t$�}|$�K�T$ QVR������L$$��t$�D$ �;M�L$w$r	�L$;M s�[��������D$ _^][��� ;]u�{ u�T$;Ur�w	�L$;M v�h �hL�h]  h��臛���D$0��_^][��� �D$][��� ����������S3�9YVu&�A��q����;�wr�A;�w�A��A�A�D$:�u�Q;Qrw�Q;r
^�Y2�[� �Q;�UWt*�q�j;�ywr�j;�w;rw��   ;z��   9YtA�q;�u(h��h��h�  h���Y賚����_]^2�[� �y;~�irw;nr
_]^�Y[� ;zw#r;js�Q�;ӉQtI��;rr�w��;rr�Q;zr(w	;jr!�d$ �Q�R;ӉQt��;rw�r��;rs�_]^[� h��h��h�  h��������_]^2�[� ����̃�(SVW�|$83�;���u9\$<t"9\$@u)h��h̟h�  h���ə����_^3�3�[��(� j�R�����uh��h̟h�  ��9\$<U�\$�\$w;��w  ��    �~ �H  �`��3�D$ wr=   w�D$    �D$ 3�j jUP�g�  �D$�F���ʉL$t"�X�x�P�@;�rw;�v+�؃�0�� �3�3ۋD$ ����;�w
r;�s����;�wZr;|$sRj jSW��  �l$��;݋�w;r;|$s3�σ�ЋÃ��9D$@r#w9L$<vj jSW�ʄ  ��;݋�r�w;|$r̓��W����W��Wj P�F�"}  �F�N��F�P �P�F�N����t�H�F�P�N�Q�@�A��N�F�F�P�H�˃������P�H�F�N�P;ʋh�~�l$(��   w;���   �X;ڋx��   w;���   ;�r&w9~r;^rw;>v�>�^�P�V�K����l$(�F+ŋ��+~�l$4�l$@�;�rw;|$<v�|$<�݋L$DWQ�N�Q�R�;�  �V��~�N^�F;�wr�;�s��F|$\$)|$<�|$D��l$@w�|$< v8�F�H�N����h��h̟h�  h��� �����]_^3�3�[��(� �D$�T$]_^[��(� ������������̃�UVW��j �t$�����l$$j jh � �͋�������u	_^]��� �F�SPQ��2��9������   W����7������   �n3ۅ�\$t~�d$ �V;ڋ�D$wmr9D$se�} tX�E�u;ƋM�}rDw;�v>+�Ƌ�L$���;�r�D$w;�v
+D$Ӌ����E�L$(PV�����tt$ߋt$�m��u��l$(����9b����u2ۊ�[_^]��� ������̸`������������S�\$V��W�~@S���l�����u ��thp�S�8����豓��_^��[� U�n<j ���[���;�t��t3hL��#�~x u5�F(;u�N,;Ou9n8t!��th�S�c8�����[���]_^��[� ]_^�   [� �����V�t$Wj j��h � @���������u_3�^� j jh � @���D$ ���������   S�GP��2��"8����tt�OQ����9����te�WR����9����tV�G,�O(PQ���7����tC�W4�G0RP���7����t0�O8Q����5����t!�W<R����5����t�GxP���3����t����`����t��tV�O@�b�����t�D$[���`����u�D$�D$_^� ��������������̋T$��8SU�l$HV3�;�W��wLr;�wF�~;���^�^�^�^��  �G���t�O ;�t	P�R����W�R�����ۋ�u��x  �F;��\  r;��@  9^�^�  9^�  ��F�P;�rFw	�H;L$Lr;�8��t�_�N�A��t�� ;�t	P�R�����VR�R����;��~u���  �F�P;�xrqw�\$L;�vkh��h��h\  h�������F�H�~�P��;�rw�>;�v��N�@    �F�V;Ћrw�V;�v�N�F_^]2�[��8� �\$L�H��t;�rw;�v+H��+�R�j Q�;w  ����n�I  h��h��hR  h���u�����_^]2�[��8� ;��  w;��  �T$L�N�F��j �U�L$4R�ΉD$4�R�������  �D$�ȅɈ\$�D$�D$   �\$uh��h̟h�  �  j��������uh��h̟h�  �n  ��$    �~ �J  ��X��3ۉD$0wr=   w�   �D$03�j jSP�}  �D$ �F���T$$t"�h�x�H�@;�rw;�v+���0�� �3�3�D$0����;�w
r;�s����;l$$w\r;|$ sTj jUW�T}  ��;l$$��w?r;|$ s7�\$�σ�ЋŃ��;�r%w9L$vj jUW�}  ��;l$$��r�w;|$ r̓��W����_O��Wj P�F�su  �F�V��F�H �H�F����t�V�P�F�P�N�Q�@�A��N�N�F�F�P�H�̓������P�H�N�V�Y;Ӌi�F�l$8��   w;���   �A;Ëy��   w;���   ;�r&w9~r;Frw;>v�>�F�Q�V�   �l$8�N+͋��+~�\$l$D��;�rw;|$v�|$��D$WP�F�P�R�x  �V��~�Nn�F;�wr�;�s��F)|$�|$�ۉ\$w�|$ v?�F�H�N�|$ �����r)�|$ ������h��h̟h�  h���_������T$,�D$(j RP���i����l$P�L$L;u;nu_^]�   [��8� _^]3�[��8� �������������Vj j ��������F    �F    ^����̃�W����ҋOu��uQQ�������G    �_��ËG����   S�XV�p;���   w;���   ;H��   r	;P��   ;Pu	;H��   +�ΉL$��L$�H��U��t�P ;�t���3ۍM QP�0M��������t\;wu��tE�ۍF �FtUSP��v  S��L�����L$��F    �G9Gu�w9Gu�w�ɉwt�q�G��P�O�H]^[�_���̃�HSVW3�W��W�t$�����\$X�D$P�L$Qh � �ˉ|$$�|$(�ih����u	_^[��H� 3��T$4R�ˉD$8�D$<�D$@�D$D�D$H�D$L�D$P�D$T�N���|$�|$$�|$(�|$ �D$ �|$��  �D$$P���"�����t  �L$ Q���~�����`  9|$U�L$8u?�����l$(�t$,�̓����;�u;�tbh$�h �h�  h���������  �W����l$(�t$,�݃����;�w'r;�s!h$�h �h�  h��裌������   ;�w;���   ;��l$0�t$4w��   v�D$0   �|$4�T$0R��J����;ǉD$��   �D$,3�3�;�re�L$(w
;�v[��L$(�|$4�t$0+��;�r
w;�v����D$�L$\PV������t/�L$Q�L$WV������D$,��;�r�w�L$(;�r�3��D$�3��D$;�t	P�J�����t$]�L$X�Z����u�D$WW�������D$_^[��H� �|$ t������W���Y���;D$ u�;T$$u	�F;D$(t�h��h �h  h���Y����D$��_^[��H� ���������j�hc�d�    PQSV�  3�P�D$d�    ��t$�����8��`/�F�d/�N�h/�V�l/3ۍN�\$�F�+���N�D$�+���^ �^(�^,�^0�^4�^8�^<�^@�^D�^H�^L�^P�^T�^X�^\�^`�^d3��Fh�Fl�Fp�^x�^y�^z�^{�^|�^}�^~�^�ƋL$d�    Y^[��������j�h��d�    PQ�  3�P�D$d�    h�   �.�����D$���D$    t��������L$d�    Y���3��L$d�    Y������������SV�������3�SS�N@�����^<�^x�`/�F�d/�N�h/�V�l/�N�F�)���N�)���^(�^,�^0�^4�^8�^<^[��������������̃�SVW�������t$ �D$P�L$Q3�h � @�Ή\$�\$ �d����u_^3�[��� �|$�\$ ��   �T$R�D$Ph � @�Ή\$�\$$��c������   2ۃ|$uz�OQ���g����tk�WR���(����t\�GP�������tM�O(Q�������t>�W0R�������t/�G8P��������t �O<Q��������t�WxR�������t����QW����t��tV�O@������t�D$ ���0W����u�D$ �D$ _^[��� ����������VW�|$��;���   SU�9���W���A���G�F�O�N�W�V�G�OQ�N�F��.���WR�N��.���G(�F(�O,�N,�W0�V0�G4�F4�O8�N8�W<�o@�^@;݉V<tj j ������3�U�ˉC�C������Gx]�Fx[_��^� ���������j�h��d�    PQVW�  3�P�D$d�    ��t$�8��D$   �d���j �~@j ���&����N�G    �G    �D$�&���N�D$ �~&�����D$����������L$d�    Y_^����������������j�h�d�    PQVW�  3�P�D$d�    ��h�   �!+�����D$���D$    t���g������3����D$����tW���M����ƋL$d�    Y_^������������VW�|$��t5h`���������t%�t$��th`���������tW�������_�^�_2�^�������������V�������D$t	V�k,������^� ����S�\$U��}V����W�   ��z����   �w��    ;}}/�E�0�Q�R�����\$����Az2ۃ�����u�_^]��[� ����   �E����   �M�@�T��R訰���\$����Azg_^2�]��[� ��tX�   ;}},��tJ�E�0�Q�R�1�����t2ۃ�����u�_^]��[� ��t�E��}�M�@�T��R�������t2�_^]��[� ������������̋D$VP��������^� ������������̋A��y3������̃�VW���w�����D$ �/  ��S�\$U������   �O�v����D$�P誯���\$����A��   �   ;���   �   �GP�(�}����\$����Au"�G�L$�R�(�_����\$����A��   ����;�|��D$][_^��� �G�v��ۍQPj j��������to���D$   ~b�   ��I �GP�(Rj j迻������u�G�Q�(Rj j褻������t �D$����;ƉD$|��D$][_^��� �D$][�D$_^��� ����������V������������^���������������W�|$��t�? tV�50!h�&��W��h�&��^_��������V�pW�x�����>�x�   p�P�:p_^����������V���F�NW�x;�v����t5�@�NWPQ�kk  �F~x~)~�F)x�v���~ u�V�V_^��VW�|$����  �w����  �L$����  � ��  �? u
� ��  �F=�  u	���|  � u����G_�����^Ã�*�V(SU�>�T$�N(�   ��  �   9F��  j j j �SQ  �G0�N�F�^�F�V��^�F�N�^�F�n������   �V�*^�F�N� ^�F�V� ^�F�N� ^�F�V� ^���   ��	�Nu�C����   }	��|3���   �V�^�F�N�^�Fq   ��  �P$�H,��҃���Ƀ�ыH��Ƀ�ыH��Ƀ�у8 �N��Ј)^�F�V�R�N�^�N�I�F�V�^�V�R�F�N�^�N�I�F�V�^���   ��	�Nu�   ����   }	��|3���   �V�^�N�F�I�V�^�F�x �Nt!�@�V�^�N�I�F�V�^�N�V�z, t�FQ�O0PQ�yO  ���G0�F     �FE   �   �N0������   9��   }���   ;�|��}���3҃�����3���ȃ~l t�� ��B��+������ˋ���+ȋ��Fq   �����~l t�O2�t����O0�k���j j j � /  ���G0�~E��   �F�x ��   �@9F �Nsn��$    �F;Fu6�V�z, t;�v+�P�F��O0PQ�yN  ���G0���,����F;F��t)�V�R�^ ��n�(�   FF �F�P9V r��F�x, t�F;�v�V+�P�G0�RP�N  ���G0�N�V ;Qu�F     �FI   �~I�   ��   �F�x ��   �V�F;Fu6�N�y, t;�v�O0+�P�F�PQ�M  ���G0���e����F;F��t!�N �^�[�͉N �N�n��u���݋F�x, t�F;�v�N+�PʋW0QR�VM  ���G0��u
�^ �F[   �~[��   �F�x$ ��   �V�F;Fu6�N�y, t;�v�O0+�P�F�PQ�M  ���G0�������F;F��t"�N �^�[$����N �N�n��u���݋F�x, t�F;�v�N+�PʋW0QR�L  ���G0��u�Fg   �~gu[�F�x, tK�N��;Nv���2����F�P;Vw5�W0�N�n�W1�F�Nj j �nj �?L  ���G0�Fq   �~ t�������� u5�F(����][_3�^Ã �\$u!;\$��t���][�G_�����^Ë\$�F=�  u� t���][�O_�����^Ã u�~t u����   =�  ��   ���   �@����SV�Ѓ���t��u�F�  ���:  ���1  ;�uW;�uV�D  ���7j j j V�D  ����u#�NL�VDf�DJ�  �FL�VD�L �Qj R�d`  ���������� �������������F����][_^Ã���   �W0�N�F�n�W1�F�N�n�W2�F�N�n�W3�F�N�n�W�F�N�n�W	�F�N�n�W
�F�N�n�W�F�N�n��O2��������O0������������F��~�؉F]3�9F[_��^Ã ����][_�F(����3�^á���G_�����^���V�t$����   �F����   W�x��*t)��Et$��It��[t��gt��qt���  t_�����^Ë@��t�N$P�F(P�у��V�BD��t�N$P�F(P�у��V�B@��t�N$P�F(P�у��V�B8��t�N$P�F(P�у��V�F(�N$RP�у�3���q��_�F    ^�����ø����^��������������̋F,�NL�VDW��F<3�f�|J��FL�VD�L �QWR�H^  ���   �@��� �����   ������   �������   �����   ���~l�~\�~t�~h�~H�V|�Fx�F`_����������̃��O|�WlSU�oxV���   �L$�O8�t$�w,�������;�v+ց�  �T$��D$    ;��   �T)��T$�)��  �T$r�l$�Wt9T$v�T$�W8�\$�8*��   �\$8\*���   �:��   �Z��:Y��   �����Y����:u_�Y����:uR�Y����:uE�Y����:u8�Y����:u+�Y����:u�Y����:u�Y����:u;�r���+ց�  ;Ս�����~;T$�Gp��},�\
��
�\$�T$�W4#ЋG@�P;D$v�l$�
����Gt;�w��^][������̋N8�FlU�l$�)��:W��  ��   �Q:P��   �����P����:u_�P����:uR�P����:uE�P����:u8�P����:u+�P����:u�P����:u�P����:u;�r�+�  ��|�Nt;��npv
_��]ø   _]��������������̃�SU�n,W��$    �~<+~t�Fl�N,+���)����;|$rc�F8U�(QP�e_  �VL�FD)np)nl��)n\�P�A���;�r+��3���f�u�N@�Սi�A���;�r+��3���f�u���|$�>� ��   �FtFl�OF8�T$��;ډD$v�څ�tM�W+ˉO�J��u��O0SPQ��%  ���u��G0SRP�cE  �G0�D$���SQP�^  ��_^t�~t��r�F8�Vl�NX���FH���J3�#FT�FH��  s��z �����_][�����QSV�t$�F���=��  W�D$��  s�D$�Ft��w�����Ft���6  Fl�N\�D$�Vl�Ft    �t;���   +ЅɉVt�Fl|�V8��3�j +�PRV��?  �Nl�>�N\�G�X�O��;�v�م�t5�P�GSRP�]  �G_X_)_�G)X���� u�O�O��z ��   �V\�Nl�F,+�-  ;��/�����|�F8��3�j QPV�G?  �Nl�>�N\�G�X�O��;�v�م�t5�P�GSRP�]  �G_X_)_�G)X���� u�O�O��z �����_^3�[YË|$��t�N\��|�F8��3�3҃���R�Vl+�RPV�>  �Fl�F\��������3�9Au����_^[����YÃ���_^[�D Y�����������SUV�t$W3ۍ�    �Ft=  s#�����Ft=  �|$s����  ����  ��rI�FH�NX�Vl�~4���N8�L3�#FT�ND�FHf�A#��V@f�z�Nl#N4�V@�J�FH�NDf�Vlf�A��t6�Fl�N,+Á�  ;�w$���   ����   ����   �Ë������F`�   �~`�O  f�Vlf+Vp�F`���  �ʋ��  f�W���  ���  ,�:��  ���� �f���  ����  ����  f�� s+���� ��,��u��   ;�u�S�������F`�p��������� �f���	  ���  3�+�9��  �����F`)Ft;��   �Ntwb��r]����F`nl�Vl�N8�D
�^H�NX��ND3�#FT�^4#ڋV@�FHf�Af�Z�Nl#N4�V@�J�FH�NDf�Vlf�A�F`�u��   Fl�Fl�N8��NX�F`    ��FH�R��3�#FT�FH�^�Fl�N8����  ���  f�Q  ���  ���  �
��  ��f���   ����   ���  3�+�9��  ���Ft���nl��������N\��|�F8��3��Vlj +�RPV��;  �Fl�>�F\�G�h�O��;�v���t5�H�WUQR�Y  �Goho)o�G)h���� u�G�G��y �	���_^]3�[ËN\��|�F8��3�3҃���R�Vl+�RPV�<;  �Fl�F\��������3�9Au����_^][����Ã���_^][�D ����QSUV�t$W�D$    �   �Ft=  s#�;����Ft=  �|$s����  ����  ��rM�FH�NX�Vl�~4���N8�L3�#FT�ND�FH�A#��V@f�z�Nl#N4�V@�J�NH�VD�D$�Flf�J�Vp�N`�Vd�T$�һ   �Nx�^`tq��;��   sg�Fl�N,+�  ;�wU���   ;�t��t���+������u;�uR�������F`�F`��w9��   t��u�Vl+Vp��   v�^`�Fx����  9F`��  f�Vlf+Vd�Fl�Nt���  �|��Fxf+��ʋ��  f�S���  ���  ,���  ���� �f���  ����  ����  f�� s���� �������� �f���	  ���  �Fx+�3�9��  ����+�Nt����Fxnl�Vl;�wN�FH�NX�n@���N8�L#V43�#FT�ND�FH�Af�DU �Nl#N4�V@�J�NH�VD�D$�Flf�J�   �Fx�u�nl�ۋFl�Fh    �F`   ������V\��|�N8��3�j +�PQV�8  �Nl�>�N\�G�X�O��;�v�م�t5�P�GSRP�[V  �G_X_)_�G)X���� u�O�O��z �>���_^]3�[YÃ~h ��   �Fl�N8�D����  ���  f�Q  ���  ���  �
��  ��f���   ����   ���  +�9��  ur�N\��|�F8��3��Vlj +�RPV�7  �Fl�>�F\�G�X�O��;�v�م�t5�H�WSQR�xU  �G_X_)_�G)X���� u�G�G�nl�Ft��y ����nl�Ft��nh�F����~h tJ�Vl�F8�D����  ���  f�J  ���  ���  ���  ��f���   ����   �Fh    �N\��|�F8��3�3҃���R�Vl+�RPV�6  �Fl�F\��������3�9Au����_^][����YÃ���_^][�D Y����������������SVW�|$3�;�ty�w;�tr9_ tm9_$th�_�_�_�G,   �F�F�F;É^}�؉F�F����Ƀ�S��q��S�NSu�:  ��  ���G0V�^(�/  ���p���_^3�[�_^�����[�̋D$3�;�U�   �  �81��  �|$$8��  W�|$;�u_�E�]�9O �Ou
�G   �O(9O$u�G$  �|$�u�D$   S�\$;�}3������~�   ���D$ ������}  �|$�r  �K����f  �|$	�[  �|$$�P  ��u�	   �W(�G Vh�  jR�Ћ������  �w�n�˽   ��^0�\$$�   �M��N4�K���NP���>�FL����FT����������F    �n,�VX�W(�G jUR�ЋN,�F8�W(�G jQR�ЋNL�F@�W(�G jQR�ЉFD�K�   ��j���  �O(�W PQ�ҋ��  ��0�~8 ��    �F�VtN�~@ tH�~D tB��t>����P�H��L$���  �T$(W���  ���   ���   �F$������^[_]��F�  ���W�G������^[_�����]�[_�����]ø����]���̋D$�L$�T$P�D$Qj jjjRP������ �����������̋T$3�;�tM�B;�tF�H�J�J�J�B0   ��H�H�H �H(�H,�H0�H8�H<��0  �@ �  �Hl�HP�HL3�ø�������̋D$W3�;���   �81��   �|$8��   V�t$;���   9~ �~u
�F   �~(9~$u�F$  �F(�N h0%  jP�у�;�u^�����_ËL$;ωF}�x�����������0�P}���Q���wV�H$�x4�������^_ËN$P�F(P�у��~^�����_ø����_�����̋D$�L$�T$PQjR�������������UV�s3�9n4W��u'�N$�S �   ���K(jPQ�҃�;ŉF4u_^�E]�9n(u�N$�   ���n0�n,�F(+{�F(;�r"�K�V4P+�QR��O  �F(��_�n0�F,^3�]�+F0��;�v��K�V4V0U+�QR�O  ��+�t"�C�N4W+�PQ�O  �V(���~0_�V,^3�]�n0�N0�F(;�u�F0    �N,;�s͉N,_^3�]���������̋T$��,��W�Y  �z���N  �z �D  �: u
�z �5  �?u�   �J�BS�_8U�*�L$�L$(����D$$�BV�w<�D$�\$�D$8�D$0    v�����^][_��,����$    �T$@�$��Z� u�   �b  ��s(����  �U ���������ڃ��D$�\$r��GtM���  uEj j j �5  �Gj�D$0�D$0�D$1��OPQ��4  3ۃ��G�D$�\$3��   ��  �G ���G    t�@0�����G��   ���������3ҹ   �����   �Ӏ���t�D$@�@���D$�  ���˃�����;O$�\$v�L$@�D$�A���V  �   ��j j j �W�  �L$L���Ӄ���	�G�A0�D$�3ۃ��\$3��  �T$@�D$�B���  ��s-��I ���P  �U ���������ڃ��D$�\$r؀��_t�L$@�A���  �� �  t�T$@�Bt��  �O ��t
��������G   t%�\$ ��j�D$$�\$%�OPQ�c3  �G�D$��3�3��   ��� s$����  �U ���������ڃ� �D$r܋O ��t�Y�G   t7�\$ �Ë�������j�T$$�D$%�L$&�\$'�GRP��2  �G�D$��3�3��   ���s$���)  �U ���������ڃ��D$r܋O ��t�Ӂ��   �Q�W �����J�G   t%�\$ ��j�D$$�\$%�OPQ�d2  �G�D$��3ۉ\$3��   �G   tn��s$����  �U ���������ڃ��D$r܋O �ɉ_@t�Y�G   t%�\$ ��j�D$$�\$%�OPQ��1  �G�D$��3ۉ\$3���O ��t�A    �   �G   ��   �O@;ȉL$v�ȉD$���   �W ��tG�R�҉T$4t<�G �@+G@�W �R�D$$�;�v+T$$�ʋT$$Q�L$8�UQ�J  �L$ �D$���G   t�D$�OPUQ�51  �L$ �G�D$��+��)O@�D$�@ �z  �G@    �   �G   ��   ���X  3��)���L$�O �ɉT$$t&�Q�҉T$4t�W@;Q s�D$4�L$$��G@�D$�|$$ t�L$;�r��G   t�T$�GRUP�0  �G�D$���L$+��|$$ �D$��  ��O ��t�A    �G@    �   �G   ��   ����  3ɍ�    �)���L$�O �ɉT$$t&�Q$�҉T$4t�W@;Q(s�D$4�L$$��G@�D$�|$$ t�L$;�r��G   t�T$�GRUP��/  �G�D$���L$+��|$$ �D$�  ��O ��t�A$    �   �G   tM��s(����  �U ���������ڃ��D$�\$r��O;�t�T$@�B`��P  3ۉ\$3��G ��t�O��	���H,�W �B0   j j j �/  �L$L�G�A0�D$���   �
  �� s/��$    ���P  �U ���������ڃ� �D$�\$r؋ˁ� �  �����3Ҋt$����ʋT$@ˉO�J03�3��
   � ��  j j j ��  �L$L�G�A0�D$���   �|$D��  � t�΃���+��   �\$�N  ��s$����  �U ���������ڃ��D$r܋˃���O�˃�����ws�$�H[���   �\$����  ���GLp��GT	   �GPp��GX   �   �\$����  ���   �\$���  �T$@�BL��   ���\$���  �΃���+�� �\$s(����  �U ���������ڃ� �D$�\$r؋Ӌ��ҁ���  ��;�t�L$@�A,��)  3ۉO@�\$3��   �O@�ɉL$��  ;�v�ȉD$�T$;�v�ʉL$���I  �T$�D$(RUP�!F  �D$ )D$)D$(D$4��)G@�D$�
  ��s$���  �U ���������ڃ��D$r܋˃�����  �ӉO`���˃������������`  �Wd�O\�\$��   ����   �Gh    �   �Oh;O\sX��s'�I ����
  �U ���������ڃ��D$r܋Wh�U��˃�f�LWp�Gh�Oh����;O\�\$r��   9Ohs �   ��Wh�U�f�DWp  Gh9Ohr捇0  �Ol��GL���  R�GTPQ�    j�GpPj �Y0  ���D$0���D$t �L$@�A��b	  �T$@�B��R	  �Gh    �   �WdW`9Wh�7  �OT�   ��OL��#Ӌ�������;։L$vD���i	  �U ����OT����ں   ��OL���D$��#Ӌ�������;։L$w�������sW������;�s*���	  �U ����L$������Ճ�;�D$r�f�T$����+�Ohf�TOp�Gh�\$�^  f�T$f���͉L$$ud�Q;�s*����  �U ����L$$����ڍQ��;�D$r���+�Oh�ɉ\$�n  �LOn�L$$�˃������L$���   f��uJ�Q;�s+����@  �U ����L$$����ڍQ��;�D$r���Ӄ����T$��������N�Q;�s1��$    ����  �U ����L$$����ڍQ��;�D$r���Ӄ����T$�������+ыL$��D$$    �WhыOdO`�\$;���   �|$ t�L$$�Wh�l$f�LWp�Gh�|$ u�OdO`9Oh������?��  ��0  �Ol��GL���  R�W`�GTPQ� 	   R�GpPj�-  �����D$0t4�L$@�D$�AЫ�  �T$@�B���  �L$@�A���  �Wl�Ol�WP���  R�GXPQ�O`�    �GdP�TOpRj�2-  �����D$0t�D$@�@���D$�;  �D$�   ��rc�|$  rY�D$@�T$�L$(�P�T$,�H�L$R�(�HP�_8�w<�(  �D$H�H�P�(�@�_8�w<���L$(�T$�D$�\$��  �OT�   ��OL��#Ӌ�������;ΉT$vD����  �U ����OT����ں   ��OL���D$��#Ӌ�������;ΉT$w�����   �����   �����L$4�ɉL$$��L$$�T$�   ��L$$��#���L$��ыOL���L$�����L$4�;�vc��    ���P  �U ����L$�������ʉT$$�   ��L$$���D$��#����L$ыOL���L$����T$$;�w��L$�T$��+��������+�L$$�����҉\$�O@u�   �i  �� t�   �Y  ��@t�T$@�B���>  ���WH�   �OH��t>;�s$���  �U ����������;wH�D$r܋OH�   ���#�W@��+��   �OX�   ��OP��#Ӌ�������;ΉT$vD���  �U ����OX����ں   ��OP���D$��#Ӌ�������;ΉT$w������   �����L$4�ɉL$$��L$$�T$�   ��L$$��#���L$��ыOP���L$�����L$4�;�v]���|  �U ����L$�������ʉT$$�   ��L$$���D$��#����L$ыOP���L$����T$$;�w��L$�T$��+��������+���@�L$$�\$t�T$@�Bh��  �������OD�WH�   �OH��tB;�s$����  �U ����������;wH�D$r܋OH�   ���#�WD��+�\$�O,+L$L$,9ODv�T$@�BH��  �   �|$ �c  �T$,+T$�OD;�v<+ʋW0;ʉL$v+ʋW4W(�L$+���W4+�W0�L$�T$$�W@;ʉT$4v����T$(+ыO@�T$$�L$4�L$�T$;�v�ʉL$+щT$�T$4+щW@�L$$��L$(��   T$$�)T$�L$(u߃@ �a  �   �V  �|$ ��  �L$(�W@����l$�L$(�   �+  � ��   �� s(���n  �U ���������ڃ� �D$�\$r؋L$,+L$�T$@JO�ɉL$,t1�W���L$(P+ȃ QRt�"  ���  �L$L�G�A0�D$��� �T$�T$,��u�� �  �����3Ҋt$��ʋ����;Ot�L$@�A0��b3ۉ\$3��   � ��   � ��   �� s+�I ����   �U ���������ڃ� �D$�\$r�;_tO�L$@�A��   ����w���^][�����_��,ËL$(�J�L$�*�B�J�w<^]�_8[�   _��,�3�3��   �D$0   ��D$0�����L$@�T$(�Q�T$�Q�)�A�( �_8�w<u�?}-�D$,;At$�D$,�\$@�j�����t�   ^][�����_��,Ët$@�l$8+n�\$,+^n^_� t4��t0� St�V�G+�RP�!  ��N�W+�QR�G  �G���F0�G�����@3Ƀ?������   �G<��F,u��t�|$Du�D$0���/���^][�����_��,ËD$0^][_��,ø����_��,Ð�EfGH�HI�I[JK�KdL�L�LM�MPN�N0O#P7S6U�U�VZWXCXY�Y�YZgM|M�M�M��������V�t$��t:�F��t3�N$��t,�@4��t
P�F(P�у��N�V(�F$QR�Ѓ��F    3�^ø����^������̋L$S�\$W��������  ��u1�D$�ʁ���  r����  �����  r����  ����_�[�V�t$��u�F^_[Ã�s?��t�ȃ������u����  r����  �q����������+��^��_�[Á��  ��   ���n^��U�������    ��  �[  ��I ���V���V���V���V���V���V���V���V���V	���V
���V���V���V���V���V��������u����q������i� ��ʸq������i� ������8���]����   ����   ��������V���V���V���V���V���V���V���V���V	���V
���V���V���V���V���V�ʃ�������r�����t�ȃ������u�q������i� ��ʸq������i� �����^��_�[���������������V���   �  3���f�0����u����	  �   f�0����u���|
  �   �d$ f�0����u����  ���  ���  ���  fǂ�   ^���Q��P  UV�t$���\  �6;ʉl$��   S}4���`  ���\  ����f;�ru��X  :�(X  w���l$���\  ����f;�r-u��(X  :�X  v+�T$���\  ��P  �L$�;�~��L$[^���\  ]YËT$[^���\  ]YÉ��\  ^]Y����������̃� �QS��I�T$�QU�)�T$$�QV�q3ɉ�<  ��@  ��D  ��H  ��L  ��P  ��T  ��X  �T$$��T  ���\  Wf�L���T  ����=  �t$�L$��  ���\  �L$�=  +���L$ �|$��t$�T$��L��L���;�~�D$��;T$$f�L�H�|$(f��H<  3�;�|��+��|$,�4��<��������  ��t�T������  �|$�D$�l$ �{����l$����   �L$�Q��T$,��H<  ���    �L$,f��H<   ��H<  u����f�: t�f��H<  ��f��H>  f���������T$��tv�t$ �I �6���t$tR���\  �M��l$��;L$$�l$,.�|�;��t�t����+�����  �l$,f��l$�t$��u��|$�t$ �����҉t$ u�_^][�� ���������̃�SU�l$VW�x3҅����D$�����J�ru��   �r��f�D�����   �����\$�D$�   ��ǋ|$�?�;�};�th;�}
f��|
  �0��t;D$tf��|
  f��
  ���
	f��
  �f��
  3҅��D$u
��   �r�;�u
�   �q���   �q��D$)\$�v���_^][����������������̃�SU�jV3���W���D$�����l$�N�~u��   �}����  �����T$�\$ �   ���    �\$��T$�;�T$$�\$�t$};��  ;���   �I ���~
  ���  �   +�;�~[���|
  ����Hf	��  ���  �P�h�H���  �P����  h�*�f��L:��T$$f���  �t$�f���|
  f��f	��  �+����  �t$�f����  ����  ;T$��   ���~
  ���  �   +�;ˉ|$~[���|
  ����Hf	��  ���  �x�9h���  �H�x����  h�*�f��L$�L�f���  �t$�f���|
  f��f	��  �|$�+����  �t$���
  ���  �   +�;ˉ|$~Z���
  ����Hf	��  ���  �x�9h���  �H�x����  h�*�f��L$�L�f���  �t$�f���
  f��f	��  �|$σ�������  ~S����Hf	��  ���  �x�9h���  �x�H����  h�*�f���򉘼  f���  �  ��f	��  ����  ��
���  �   ��   ���
  +�;ˉ|$~Z���
  ����Hf	��  ���  �x�9h���  �H�x����  h�*�f��L$�L�f���  �t$�f���
  f��f	��  �|$σ�������  ~S����Hf	��  ���  �x�9h���  �x�H����  h�*�f���󉘼  f���  �  ��f	��  ����   ���
  +�;ˉ|$~Z���
  ����Hf	��  ���  �x�9h���  �H�x����  h�*�f��L$�L�f���  �t$�f���
  f��f	��  �|$σ����	���  ~P����Hf	��  ���  �x�9h���  �x�H����  h�*�f�������  f���  ���f	��  �����  �L$3��ɉT$u
��   �~�;�u
�   �y���   �y��D$)l$ �M���_^][��������Q���  ��S�\$UVW�   ~^�t$����������Hf	��  ���  �P�h���  �H�P����  h�\$ �*�f�������  f���  ��T$��������f	��  �����  ���  ��~_�t$�������H�\$f	��  ���  �P�h���  �H�P����  h�\$�*�f�������  f���  ��T$�����f	��  �����  ���  ��~[�s�����H�\$f	��  ���  �P�h���  �H�P����  h�\$�*�f���􉐼  f���  ��S���f	��  �����  3�����   ��I ���  ����L�~\���~
  ����Hf	��  ���  �P�h���  �H�P����  h�\$ �*�f���󉐼  f���  �f���~
  f��f	��  �����  �;��m����L$������   �����L$_^]������	  [�������̃�S�\$U3�9��  VW�9  ��$    ���  �,J���  �4����L$���  ��   �|��   +�;�~\�4�����H�\$f	��  ���  �P��@���  �H�P����  �@�\$�*�f��L:�f���  �  f��f��f	��  ��r  �� ����  �   +�;ˉ|$�|$ �T$~c���  ����Hf	��  ���  �P��@�H���  �P����  �@�*�f��L$�T
����  �T$f���  �f���  f��f	��  �|$ω��  �<�ج���\$ tz+4� ����  �   +�;�~Q����Hf	��  ���  �P��@���  �H�P����  �@�\$ �*�f��L:�f���  ���f	��  ω��  ����   s	�� �������� ��L$$�T����  �   +�;ΉT$~c�T$$�4�����Hf	��  ���  �P��@���  �H�P����  �@�\$ �*�f��L$�T
����  f���  ��t$$f�4�f��f	��  ʉ��  �4�`����~   ���  +,����   +�;�~U����H�\$f	��  ���  �P��@���  �H�P����  �@�\$�*�f��L2�f���  ���f	��  Ή��  �L$;��  �������  ���  �   +�;�~s��   ����H�\$ f	��  �P���  ��@�h�H���  �\$ �)���  �@�*�f��L:�_���  f���  ��  ^]���  [���f��   f��f	��  �_���  ��  ^]���  [��������3����   f�9 u������	|��	��   �   ���   �I f�y� ��   f�9 u5f�y u?f�y uIf�y uSf�y u]������ |ȋ3Ƀ� ���J,Ë3Ƀ��� ���J,Ë3Ƀ��� ���J,Ë3Ƀ��� ���J,Ë3Ƀ��� ���J,Ã��3Ƀ� ���J,�����̋��  ��Su9���  �P�H��@���  �H�P��@3ɉ��  f���  [Ã�|)�H�P���  �f���  �@���  �f���  [�����������̋��  ��SV~=���  �P�H����  �P�   p�H�p3�^f���  ���  [�3�;�~�p�P���  �2�@^f���  ���  [��������������SVW�ً��t����|$ ǀ�     �   t:�H�P�x�H�P�<x�PU�h���ш*x�h�P���ш,*x]��t�H�P+߉\$���\$x���u�_^[��������������̋T$���   ��  ��|
  ��0  3����	  ǂ   ���$  ǂ,  �ǂ8  �f���  ���  ǂ�     �l��������������̃� V�t$3ɸ   +֍4Bf�t4f�f���f�LD����~�3���|<U�T���t*�DT�ȃ�f�DT3����Ń���������f����;�~�]^�� ����������̃��D$SUW�8�@�H�(3҃��3�;ʉL$�\$��P  ǆT  =  ~7f9�t#��P  ��P  ���\  �D$��0X  ���f�T���;D$|Ƀ�P  }R��}�����3���P  ��P  ���\  f�� ��X  ���  �;�t�D�)��  ��P  |��\$�L$�Y��P  �+�����|U���f���������}�\$��$    ��P  ���\  ��`  �����P  j�Ɖ�`  �%�����`  ����T  ��T  ���\  �T  ��T  ���\  f��f���f����X  ��.X  :�r����ɀ���X  ��f�L�f�L���`  j�ƃ���������P  �D�����T  ���T  ��`  �L$���\  ���?����\$��<  ����_][������������V����  ���   V�+�����(  ���	  V������0  P��������   ��I ��L�f���~
   uk��K�f���~
   u8��J�f���~
   u5��I�f���~
   u2����}��L@��  ^Ã��L@��  ^Ã��L@��  ^Ã��L@��  ^�������̋D$���  ��~iSV�t$����Hf	��  ���  �P����  �@�H�P����  �@�*�f��L$��󉐼  �T$f���  ^[j�:���YËT$������  �L$f	��  �T$j����Y�̋D$���  �   ��SVWf	��  ���   ~J���  �P�H�p���  �H�P����  p�*ʿ   f���󉐼  f���  �	�����  ���  3���f	��  ��	~G���  �P�H�p���  �H�P����  p�*�3�f�������  f���  �	�����  �-������  ���  +у���	��   �   ��f	��  ��~J���  �P�H�p���  �H�P����  p�*ʿ   f���󉐼  f���  �	�����  ���  3���f	��  ��	~X���  �P�H�p���  �H�P����  p�*�3�f�������  f���  �M���_^ǀ�     [Ã����  �1���_^ǀ�     [����QS�\$V�t$���    W�D$    ~W��v��x,u��� �����  Q�d�����$  R�X��������N������  ���  ��
��
����;ʉD$w��K�эC;�w�D$��t�|$ WSPV��������U  ���   ��   ;���   ���  ���|$ �W~R�����Nf	��  ���  �F��F���  �N�F����  �F�*�f���󉞼  f���  ���f	��  �����  �D$��(  ��  ��P��Q��R���������	  P���   Q����������   ���  ���|$ �G~R����Nf	��  ���  �V��F���  �N�V����  �F�*�f���󉖼  f���  ���f	��  �����  h��h(����Q�������������_t��^[������^[Y���V�����t)��$    ��t�3Ё��   ��3������uރ� SW��  ����3�������܁��   ���3����%�   ��3����3����3Q�������%�   �����3���ځ��   ��3����3����3A������܁��   ���3����%�   ��3��3��3Q����%�   �����3���ځ��   ��3��3��3A������܁��   ���3����%�   ��3��3��3Q�����%�   �����3������3�����   3��3�������܁��   ���3����%�   ��3����3���� 3Q�����%�   �����3������3�����   3�����&�����rH����3���������   �<����3<������3<��%�   3<��������u���_[t��3Ё��   ��3������u���^���������������̋L$��u3�ËT$�D$�H����������̃�<SUVW�L$P�A�Q�X8�)���T*��T$�q�I��+T$T��֍�1�����T$8�P(�L$,�H,�T$(�P0�L$<�H4�T$D�PL�L$@�HP�T$ �L$$�HT�   ��HX�D$�x<�D$T   �D$T�����l$�T$H���D$0���s$�E��������������E ���l$؃��L$ #Ӌ�����������+���tC��uK��@�G  �   �L$T�ʋT$T������#�ЋD$ ������������+���u�������`  �����D$Tt.;�s�E�������l$؃��ʸ   ����#�D$T��+���s$�U���E�σ��������ډl$؃��L$0�T$$#ˋ�����������+���T$u?�d$ �@�e  ���D$�   ��L$$��#�Ћ�����������+���T$t�����;��T$s,�U��������l$�;�s�U������l$ڃ��   �ы���+���#ӋʋT$ыȋ�+D$8��;ЉT$�O  ��+�;l$<��  �L$@�D$D������L$4u,�D$(+��;l$T��   )l$T�d$ �A�������u��t;�sR��+�T$(+��;l$Tsb)l$T�d$ �Q�������u�;D$T�L$4s@)D$T��A�������u���+L$�"+��;l$Ts)l$T�A�������u���+ʋD$T��v>�P�������������A�l$T������Q������A�������uӋl$T��t�Q�������v�A����l$�T$;���   ;t$,��   �T$H�������+����    �H���N�P��������H������L$T�����L$Tw̅�t��P�������v��@���냋L$P�T$�l$�AH��   �3�D$P�@h���� t�T$�   ��D$P�@���L$�   �T$����+����+��ϸ   ���L$P+Ճ���#؍E��F�A�D$,+�  �A�D$�Q�x<_^]�X8[��<��������̃�|��$�   3���SU��$�   V�D$H�D$L�D$P�D$T�D$X�D$\�D$`�D$dv��    �LE f�DLH�LLH��;�rꋴ$�   ��D$�   f�|\H u����s�;É\$v�\$��u7��$�   �f�\$�D$@�D$�L$�
� ��
� �   ^]3�[��|þ   f�|tH u<f�|tJ u"f�|tL uf�|tN uf�|tP u����v�������������9t$s�t$�   ��$    �LDH�+�x(����v��W��$�   ~��t��t_^]���[��|�^]���[��|�f�D$n  �   ��$    f�LlfLL����f�Llr鋜$�   3���v3f�|E  t$�TE �LTl��$�   f�J�TE f�DTl�TTl��;�r͋ǃ� �����t=��t�D$4h��D$0���T$,�9���-  �D$4�(�-  �D$,   ���$�   �D$4�D$,   �D$0��$�   ��L$ �L$�   ���T$83�3ۃ��P��t$�D$<�D$(�T$@u=�  �o  ��$�   �D$$�L$�t$$��T$,*ˈL$��;�}�D$ f�D$�-~��T$0���T$4f��L$f�D$��D$`f�D$  �L$�D$<+˺   ��ˋ���L$ �D$D�4�    ����|$��$    +�+΅��9u��T$�J��   ����t
�d$ ���u���t�H�#�ȋ��3�f�DTL���DTL�D$$f��u ;T$��   �T$$���$�   �A�T$;T$������t$@#�;t$8�t$H�������u�\$�D$ �L$D���L$+ˉT$ �   ���;T$s&�tTL�d$ �>+ǅ�~�������;T$r�t$H�   ��D$(��$�   �D$<u�|$(�  ��   �֋�$�   �����D$�D���L$ +����T$8f�L��?�����$�   ��*Å��D$@�D$f�D$  t`�t$ ��$    ��t�L$@#�;L$8t�D$�73ۉD$�D$�Ћˋ���L$���J��   ����t	�I ���u���t�H�#�ȋ�u��T$(��$�   ��    �T$_^]�3�[��|�_^]�   [��|�jD�.��X  h���M��!-���e� �E�P�M��a,��h��E�P�E��&��
  �jD�Q���W  h���M���,���e� �E�P�M��",��h8%�E�P�E��(�
  �U��QQSV��3�9E��M��   t	�U�E�;�t��C��E��>"u3�9E��E�"��F�E��4���t��C��E���PF�[  ��Yt���t��CF�}� �Mt4�}� u��}� t�}�	u���t�C� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E����t��C�3�B3��FA�>\t��>"u3��u�}� t�F�8"u���3�3�9E����E����I��t�\C���u���tA9M�u< t8<	t4��t*��P�-Z  ��Yt��t��CF���C���tF��F�o�����t� C��M�����E��^[t�  ���U��QQSVW3�9=��u�d  h  �H�VW�L� �� ���;ǉ5��t�8 ��u�ލE�PW�}�3��������E�=���?YYsO�M����sG�����;�r;P��\  ����Yt.�E�P�7V�}���������E�YHY����5����[  �������_^[��Q���#d  Y�V��������D$tV�O���Y��^� �D$��	Q��	P�gd  ��Y�Y@� U��QS�E���E�d�    �d�    �E�]�m��c���[�� XY�$��U��QQSVWd�5    �u��E���j �u�u��u�_� �E�@����M�Ad�=    �]��;d�    _^[�� U���SVW��E�3�PPP�u��u�u�u�u��o  �� �E�_^[�E���]�V��t$�N3���  j V�v�vj �t$$�v�t$$�o  �� ^�U���8S�}#  u�ˉ�M�3�@�   �e� �E����  �M�3��E��E�E�E�E�E�E�E �E��e� �e� �e� �e�m�d�    �E؍E�d�    �E�   �E�E̋E�E���r  ���   �EԍE�P�E�0�U�YY�e� �}� td�    ��]؉d�    �	�E�d�    �E�[��U��QS��E�H3M��  �E�@��ft�E�@$   3�@�l�jj�E�p�E�p�E�pj �u�E�p�u�pn  �� �E�x$ u�u�u����j j j j j �E�Ph#  �������E��]�c�k ��3�@[��U��QSVW�}�G�w�E����-���u�^u  �M�N��k���M9H};H~���u	�M�]�u�} }ʋEF�0�E�;_w;�v�u  ��k�E�_^[�ËD$V�t$��q  ���   �F�|q  ���   ��^��mq  ���   ��;L$t	�@��u�@�3��V�Kq  �t$;��   u�:q  �N���   ^��*q  ���   �	�H;�t���x u�^�t  �N�H^�U����  �e� �M�3��M�E��E�E�E@�E���M��E�d�    �E�E�d�    �uQ�u�ut  �ȋE�d�    ����;  u���t  ���` �` � ��S�\$VW�������t&P�P  ��FV�  ��YY�Gt�3VP�`u  ����g �G   ��_^[� S�\$V�����C�F���CWt1��t'P�2P  ��GW�?  ��YY�Ft�sWP�u  ���	�f ��F_��^[� �y ��t	�q��  YËA��u�$��V��������D$tV�h���Y��^� ����&��&���&\��&���&��&��&��&��&���&�������  �|$ �T�t�h  �����̃��$蝂  �   ��ÍT$�H�  R��<$�D$tQf�<$t� �  �   �u���=P� �s�  �   �@ �p�  �  �u,��� u%�|$ u���Ձ  �"��� u�|$ u�%   �t����-�&�   �=P� ��  �   �@ ��  Z�U��V�uW3�;�u3��e9}u��  j^�0WWWWW�  �����E9}t9urV�u�u�.  �����uW�u�  ��9}t�9us�  j"Y����jX_^]�U��EVW3�;�tG9}u蚂  j^�0WWWWW�:  �����)9}t�9Es�u�  j"Y�����P�u�u�  ��3�_^]ËD$�X��U��$X�����(  �  3ŉ��  V���   ���   ���   �]|�ux�}tf���   f���   f�]pf�Elf�ehf�md����   ���  ���  ���   �E�  ���   �@�jP���   �E�j P��   �E��EЍE؃��E�  ��u��E��$ j ���  �E�P� ��u��uj辁  Yh  �� P� ���  3�^������Ũ  ��U���5X��aj  ��Yt]��j�x�  Y]�����3�PPPPP��������U��� �EVWjY�D��}��E��E��_�E�^t� t�E� @��E�P�u��u��u��( �� �����������̋T$�L$��ti3��D$��u��   r�=�� t�>�  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�������U��WV�u�M�}�����;�v;���  ��   r�=�� tWV����;�^_u^_]�́  ��   u������r*��$�����Ǻ   ��r����$����$�����$�(������#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ���������r���$����I ��x�p�h�`�X�P�H��D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�����������̒�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�0������$����I �Ǻ   ��r��+��$�4��$�0��D�h����F#шG��������r�����$�0��I �F#шG�F���G������r�����$�0���F#шG�F�G�F���G�������V�������$�0��I ���������'��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�0���@�H�X�l��E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_���5L���e  ��Yt��j芀  jj �c�  ���h  �U��WV�u�M�}�����;�v;���  ��   r�=�� tWV����;�^_u^_]�=~  ��   u������r*��$�$���Ǻ   ��r����$�8��$�4���$����H�t���#ъ��F�G�F���G������r���$�$��I #ъ��F���G������r���$�$��#ъ���������r���$�$��I �� �������ؕ�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�$���4�<�H�\��E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��������$�p��I �Ǻ   ��r��+��$�Ė�$����Ԗ�� ��F#шG��������r�����$����I �F#шG�F���G������r�����$�����F#шG�F�G�F���G�������V�������$����I t�|��������������D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�����Зؗ����E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� �����������̃=�� t-U�������$�,$�Ã=�� t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$�������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uZ�}  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�U}  �����$�T$�D$�   ��ÍT$�v  ��P��<$f�<$t��u  ��  ��T$��  ���   ��u  ��   �  ���   �L$���S  ���ou  ��u���=P� ��u  �X �   �4v  �=P� ��u  �X �   ��t  ZÍT$�hu  �D$uA�3���   ���D$u����   �3��3�%�� D$uÍT$�+u  �D$��%  ����� =  �uT$u���u���t��Q���$�\$��q��  ��Y�a���t���5u  �   �B����D$%�� D$������؋D$%���D$t=�f   �l$���D$�   t�- )��t��   ����������t  ����t  ������t  ���   ��������������-�&�   ���������ٱ ����u�P �������ٛ���u������U��� S3�9]u�u  SSSSS�    �)���������M�E;�t�V�E�E��EPS�u�E�P�E�����E�B   �W�  ���M��x�E����E�PS�܉  YY��^[�ÍD$Pj �t$�t$�t$�z�  ���U��Q�E��SVW�  �@ ��   Wj ��P�< ����u3��  V�>�8 ��Vj u��P�4 �ދF�~�E�F�E�F�E����  ��P�4 �E��t�� �  �M��x��E�����j����������=|�臚  ��Y�s���� a  ��u
�ʚ  �`����Ù  �0 ����~�  �`���  ��}��]  ���r����| 耗  ��|j �\A  ��Yu�\��   ��  ��3�;�u59=\�������\�9=��u�B  9}u{��  �o]  �2�  �j��uY�,]  h  j��F  ��;�YY�����V�5�&�5���\  Y�Ѕ�tWV�c]  YY�, �N���V�{  Y�m�����uW�_  Y3�@_^[�� jh��螛  ����]3�@�E��u9\���   �e� ;�t��u.�d���tWVS�ЉE�}� ��   WVS������E����   WVS�:+���E��u$��u WPS�&+��Wj S�����d���tWj S�Ѕ�t��u&WVS�~�����u!E�}� t�d���tWVS�ЉE��E������E���E��	PQ讚  YYËe��E�����3����  Ã|$u蚜  �t$�L$�T$�����Y� QSUVW�5���$[  �5�����t$�[  ��;�YY��   ��+ލk��rxV��  ��;�YsJ�   ;�s���;�rP�t$�cE  ��YYu�F;�rCP�t$�LE  ��YYt3��P�<��3Z  Y����t$�$Z  ���W�Z  Y����D$Y�3�_^][Y�Vjj �D  ��V��Y  ����������ujX^Ã& 3�^�jh��蟙  ��=  �e� �u�����Y�E��E������	   �E�軙  ��=  ��t$���������YH�jh ��Q�  �e� �u;5P�w"j�7�  Y�e� V�y�  Y�E��E������	   �E��]�  �j�4�  Y�U�l$�����   S�< VW3�95T���u��u  j�#t  h�   ��<  YY�`���u;�t���3�@P���uU�S���;�Yu;�u3�G�����WV�5T��Ӌ���u&9��j_tU賧  ��Yu����o  �8��o  �8_��^[]�U葧  Y��o  �    3�]�jh ��?�  �u��tu�=`�uCj�$�  Y�e� V蒜  Y�E��t	VP讜  YY�E������   �}� u7�u�
j��  Y�Vj �5T��4 ��u�Wo  ���D P�o  �Y��  ���������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU��  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u镦  ���$�rm  �   ��ÍT$�m  R��<$tmf�<$t��l  =  �?s+��������������=P� �@m  �   �` �=m  w:�D$��%�� D$u)��   ����-�&t�����l  ���� u�|$ u����-�&�   �=P� ��l  �   �` ��k  Z����������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU��  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�Ū  ���$�"l  �   ��ÍT$��k  R��<$tmf�<$t�k  =  �?s-����������������=P� ��k  �   �p ��k  w8�D$��%�� D$u'��   ���t��������Bk  ���� u�|$ u����-�&�   �=P� ��k  �   �p �j  Z����������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�)�  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�ծ  ���$��j  �   ��ÍT$�}j  R��<$tPf�<$t�-H�������z�=P� ��j  �   �� �j  �-J���������z��������j  ���� u�|$ u����-�&�   �=P� �Wj  �   �� �`i  Z�������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU驯  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�U�  ���$�i  �   ��ÍT$�Mi  R��<$tPf�<$t�-H�������z�=P� �|i  �   �� �yi  �-J���������z���������h  ���� u�|$ u����-�&�   �=P� �'i  �   �� �0h  Z�������̃=�� ��  ���\$�D$%�  =�  u�<$f�$f��f���d$�ڲ  � �~D$f(��f(�f(�fs�4f~�fT��f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$讯  ���D$��~D$f��f(�f��=�  |!=2  �fTp��\�f�L$�D$����f���fV��fT��f�\$�D$���������������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU陲  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u�E�  ���$�Bg  �   ��ÍT$��f  R��<$t6f�<$t�-H�����=P� � g  �   �� �g  �f  �&��� u�|$ u����-�&�   �t���뻸   �=P� ��f  �   �� ��e  Z������̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�i�  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u��  ���$�"f  �   ��ÍT$��e  R��<$tL�D$f�<$t�-H��  �t^�   �uA������=P� ��e  �� �   ��e  �   �u�ԩ�� u�|$ u%   �t����-�&�   �"�8e  ���� uŃ|$ u����-*)�   �=P� ��e  �� �   �d  Zú� �!�  �� 霵  �Ƀ=T�t�����  �����z����U��E�MV�p��uW3��;ωMu ;�t�?f  WWWWW�    �������3��9}v�9}t�;�Sv	3�[_^]�3�����tK�E�e��u�C��EE��W�u�U��YYt#}+}�} ��u�C��
�E��}��9uv�몋��;�t��u�u�U���Y��#EY��������������̋L$W����   �|$V��   St�����t9��   u�����~Ѓ��3�� �t�G���t!��t�  � t�   �uσ�����������t$��   u	����u\�"�����t=�����t)��   u����u8�˃�t��������t��u�[^�D$_È�D$[^_É����tȺ���~�Ѓ��3��� �t܄�t΄�t*��  � t��   �uĉ�D$[^_�f�3ҋD$�W[^_�f��D$[^_�����������̋L$W����   VS�ًt$��   �|$u����   �'��������t+��t/��   u����ua��t��������t7��u�D$[^_���   t�������   ��   u����ut�����u�[^�D$_É����t�����~�Ѓ��3��� �t܄�t,��t��  � t��   �uĉ�����  �����   ��3҉��3���t3������u����w����D$[^_������������̋L$WSV��|$��to�q��tU���L$���:�t��t���:�t
��u�^[_3�Ê��:�u�~��a��t(���:�u��A��t�f���:�t��3�^[_�����  �G�^[_Ë�^[_ËD$��V���F uc��M  �F�Hl��Hh�N�;�-t��,�Hpu���  ��F;`%t�F��,�Hpu�L8  �F�F�@pu�Hp�F�
���@�F��^� �D$V3�;�u�b  VVVVV�    ���������^Ë@^�U����MS�]VW3�9}�M��]�t!9}t;�u��a  WWWW�    W�g�����3�_^[�Ëu;�t���3��u9Ev!���tSWQ�������;�t����3��u9Ew��}�}f�F�}���t�F�E���E�   ����   f�FtD�F��t=�5  ;؋�r��;}���   W�6�u��u������)~>}�+߃�)}��}��   ;]�rh�}� t����3�;�v	���u������u��+������;�w��;E���   P�u�V����YP���  ������   �����   E�+�)E��(V���  ���Y��   �}� tN�M��E���FK�M��E�������E����3��}�t�uV�u�������A`  VVVV� "   V�t����}�t�uj �u�W������`  � "   3�PPPPP�G����N ��+�3��u�?����N��jh@��]�  3��u�9ut79ut29uu5�}�t�uV�u��������_  �    VVVVV�Q�����3��Z�  ��u��  Y�u��u�u�u�u�u�������E��E������   �E����u���  Y��t$�t$�t$j��t$�S������U��Q�e� S�]��u3��   ��Wru�{���vn�M�E�������tR:Q�uM�P���t<:Q�u7�P���t&:Q�u!�P���t:Q�u�E�9}�r��?�@��I��F�@��I��<�@��I��2�@��I��(�M�E����t:u@A�E�9]�r�3�_[��� �	+���jh`���  �M3�;�v.j�X3���;E�@u�T^  �    WWWWW�������3���   �M��u;�u3�F3ۉ]���wi�=`�uK������u�E;P�w7j�u�  Y�}��u趒  Y�E��E������_   �]�;�t�uWS������;�uaVj�5T��< ��;�uL9=��t3V�X�  Y���r����E;��P����    �E���3��uj��  Y�;�u�E;�t�    ���"�  �U��Q�e� W�E�P�u�u�����������uV�u���t�1]  ��t�(]  �0^��_��jh��葅  �]��u�u�t���Y��  �u��uS�$���Y�  �=`���  3��}�����  j�C�  Y�}�S貉  Y�E�;���   ;5P�wIVSP苎  ����t�]��5V�X�  Y�E�;�t'�C�H;�r��PS�u�����S�b�  �E�SP胉  ��9}�uH;�u3�F�u������uVW�5T��< �E�;�t �C�H;�r��PS�u��k���S�u��6�  ���E������.   �}� u1��uF������uVSj �5T��P ����u�]j�v�  YË}����   9=��t,V�m�  Y��������[  9}�ul���D P�^[  Y��_����   �[  9}�th�    �q��uFVSj �5T��P ����uV9��t4V��  Y��t���v�V���  Y�;[  �    3����  ��([  �|�����u�[  ���D P��Z  �Y����jh���v�  3��]3�;���;�u��Z  �    WWWWW����������S�=`�u8j�5�  Y�}�S複  Y�E�;�t�s���	�u���u��E������%   9}�uSW�5T��T �����6�  �3��]�u�j��  Y�����������̺`1��  �`1�\�  jh��贂  �e� �Mx:�M+M�M�U��E�E�E� �E��E��8csm�t�E�    �E���WH  �e��E�����誂  � jh���V�  �e� �u���EE�e� �Mx)u�M�U���E�   �E������   �_�  � �}� u�u�u�u�u�@����jh ���  3��E��E��E�E�;E}�u���Uu�u�E����E�   �E������   ���  � �}� u�u�u��u�u������������Q�L$+ȃ����Y����Q�L$+ȃ����Y�������̃=�� tn���\$�D$%�  =�  u�<$f�$f��f���d$uA�-�  ��=�� t<���\$�D$%�  =�  u�<$f�$f��f���d$u���  �Z)鐩  �Z)鳧  ����̃=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�Y�  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u��  ���$�V  �   ��ÍT$�=V  R��<$tTf�<$t�-H������z�؃=P� �jV  �    �!�gV  �-J���������z�����������U  ���� u�|$ u����-�&�   �=P� �V  �    �!�U  Z�jh ��  3ۉ]�3��};���;�u�W  �    SSSSS������3��y3��u;���;�t�3�8��;�t��}�  �E;�u��V  �    �ʉ]�8u �V  �    j��E�Ph  �x�  ���P�uVW��  ���E��E������	   �E��3  ��u���  Y�VW�|$3�;�u�UV  j_VVVVV�8����������&h�   �t$�t$������;Ɖt3���V  � _^�SV�t$W3����;�u�V  WWWWW�    ��������B�F�t7V�  V����  V����P�.�  ����}�����F;�t
P�����Y�~�~��_^[�jh@��~  �M��3��u3�;���;�u�U  �    WWWWW�����������F@t�~�E��~  �V�]�  Y�}�V�/���Y�E��E������   �ՋuV��  Y�U��$X����(  �����  3ŉ��  SV���  WV�������3�9FY�}�}�FjPPW���  �ڃ��ۉE��]�|��s
�����]  �ǃ�k�8�������E�� ǊH$���f�F�M�u�F�M��+�ڋ����  ��^��+Ӌ^���U��  �}���   3�9X0��   ��9^�U�u�E��U���  S�p,�p(�u���  ���E�� ���;w(�U��N���;W,�E���S�E�Ph   �E�P�7�X ���'���S�u��u��u����  ��;�����;������M��}�;������;��E�t4�T�O;�s+���u�J�;�s�H�9
u��������-�@;�uЍM�+�3��U��  �@�t�V�	�:
u�E�B;�r�U�U�u�E���   ��x��CS  �    �m����V����   �V��u!U��   +N��@�����   jj j �u����  ��;E�u ;U�u�F���8
uC@;�r�f�F  �Lj �u��u��u���  �����������������   ;�w�N��t	f�� ��t�^�E�� �D8tC�}�u��)]��]� �}�u�m��E�3�E�U����  _^3�[������Ũ  ��jh`��z  �u�F�  Y�e� �u����Y�E��U��E������   �E��U���z  ��u�|�  Y�U���SVW3�9}t$9}t�u;�u��Q  WWWWW�    ������3�_^[�ËM;�tڃ��3��u9Ew͋}�}f�F�M��}��t�F�E���E�   ����   �N��  t/�F��t(��   ;؋�r��W�u��6����)~>��+�}��O;]�rO��tV�  ��Yu}�}� ��t	3ҋ��u�+�W�u�V�����YP���  �����ta;ǋ�w��M�+�;�rP�}��)�E�� VP�e  ���YYt)�E��FK���E��E�   ���A����E������N ��+�3��u������N �E���jh���y  3�9ut)9ut$3�9u��;�u �zP  �    VVVVV������3��"y  ��u�e�  Y�u��u�u�u�u�@������E��E������   �E����u��  Y�SV�t$�F�Ȁ�3ۀ�u?f�t9�FW�>+���~,WPV�����YP��  ��;�u�F��y����F��N ���_�F�f �^��[�V�t$��u	V�3   Y^�V������Yt���^�f�F @tV�p���P�$�  YY���^�3�^�jh����w  3��}�}�j��{  Y�}�3��u�;5@���   �,���98t^� �@�tVPV�|�  YY3�B�U��,����H���t/9UuP�P���Y���t�E��9}u��tP�5���Y���u	E܉}��   F�3��u�,��4�V�{�  YY��E������   �}�E�t�E��ow  �j�Fz  Y�j����Y�U���S3�9]VW��   �u�M������9]u.�qN  SSSSS�    ������8]�t�E��`p������   �};�t˾���9uv(�2N  SSSSS�    �������8]�t�E��`p����`�E�9Xu�uW�u��  ��8]�tD�M��ap��;�E� �M�QP��  �E����M�QP��  ��G�Mt;�t;�t�+����3�_^[��U��V3�95��u99uu�M  VVVVV�    �1����������'9ut܁}���w�^]���  V�u�u�u������^]�U��V�u�F��u�;M  �    ����f���}�FuV�V�  E�e YV������F��Yy����F��t�tf� u�F   �u�uV�����YP�4�  3Ƀ������I��^]�jh���8u  3�3�9u��;�u�L  �    VVVVV�G���������>�};�t
��t��u��u��  Y�u�W�u�u�������E��E������	   �E��u  ��u��  YËD$V3�;�u�2L  VVVVV�    �������3�^Ë@��^�������������SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� �T$V�t$W��H�F��w�� �
�y�B��w�� ��t;�t�_+�^�U���S�u�M�����3�9]u.�LK  SSSSS�    �������8]�t�E��`p������   W�};�u+�K  SSSSS�    ������8]�t�E��`p������U�E�9XuW�u�@���YY�4V�E� �M�QP��   �E����M�QP��   ��G;�t;�t�+���^8]�t�M��ap�_[��U��V3�95��u09uu�J  VVVVV�    �����������9ut�^]����V�u�u�������^]ËD$��t���8��  uP�`���Y������U��WV�}�׋�3�������t��;�s�&���'�������^_��U���SV�u�M��>����]�   ;�sT�M胹�   ~�E�PjS��  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�<�  ��YYt�Ej�E��]��E� Y��=I  � *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P謯  ��$���o�����u�E���M�3��e���}� t�M��ap�^[�Ã=�� u�D$�H���w�� �j �t$�����YY�U���SV�u�M�� ����]3�;�u/�H  VVVVV�    �2������}� t�E��`p�������   W�};�u/�\H  VVVVV�    ��������}� t�E��`p������   �E�9pu:�f=A r	f=Z w�� ���f=A r	f=Z w�� CCGGf����t8f;�t��1��M�QP菳  ����M�QCPC�}�  ��GGf����tf;�t�����+��}� t�M��ap�_^[��V3�95��Wuq�|$;�u�G  VVVVV�    �+����������[�T$;�t��f=A r	f=Z w�� ���f=A r	f=Z w�� GGBBf;���tf;�t�����+��V�t$�t$�f�����_^�U��� S3�9]u �G  SSSSS�    ����������   �M;�V�ut!;�u��F  SSSSS�    �q���������S����;ȉE�w�M�W�u�E��u�E�B   �u�u�P�u��\  ��;��t�M�x�E����E�PS�[  YY��_^[���t$j �t$�t$�t$�8������U��� S3�9]u �5F  SSSSS�    �����������   �E;�V�ut!;�u�F  SSSSS�    ����������t=���?�E�B   �u�u�v	�E�������E�W�u�E��u�uP�"�  ��;��t5�M�x
�E���E���E�PS�IZ  YY�M�x�E����E�PS�1Z  YY��_^[���t$j �t$�t$�t$�������jh����m  3ۉ]�j�q  Y�]�j_�}�;=@�}W�����,��9tD� �@�tP�o���Y���t�E��|(�,���� P�\ �,��4����Y�,��G��E������	   �E��m  �j�_p  Y�jh��-m  3�3�9u��;�u�D  �    VVVVV�<���������_跸  j [�Pj轹  YY�u�蠸  �P���  Y���EPV�u舸  �P�[Z  �E��x�  �PW�G�  ���E������	   �E���l  ��R�  �� Pj边  YYá  ��3�9p������jh(��hl  3�3�9]��;�u ��C  �    SSSSS�w����������   3��u;���;�t��F@��   V����Y���t.V�t���Y���t"V�h������<���V�X���YY��k�8���)�@$u�V�;���Y���t.V�/���Y���t"V�#������<���V����YY��k�8���)�@$��:����u�h  �E�V��  YY�]�V�t�  ��V�u�j�u������E�VW���  ���E������   3��M�9M���H�k  ËuV�/�  Y�U���V�uW3�;��}�u�B  j^WWWWW�0�<��������  j$h�   V�����E��;�tˋ�@;ǉM��E�|;�s�RB  j^�0����|
����o@�w�SWh�3�PQ�w�  �ȃ�F��+  ���  ���y�jd�}��M�؋Ǚ_��j�h����+؋E��������D��A��ڙRP����+��j ��Q SRP�����}��U�}� M|��sG�E��ǀ3��U� �ȁ�  ��EyI���Aujd�Y����u�El  ���  ����uA��U� �2�E�ȁ�  �yI���Au
jd�Y����u�El  ���  ����u�E�   �Ej S�u�FW�o�  j��F�h����RP������U�}� ��1u��1�F3�A9B}��A9�|���Q I�N+�j �F�ES�p�0��  j��Y���3�Sh  �u�W�V���  j��F�h����RP�W���S�U�j<�u�W���  �Fk�<+��^ �>3�[_^��V�f�  ����u^��t$V�������Y��Y#�^�U��QQ�E�P�` �E��M�j  ��*h��� ��!Nb�QP� ����M��t��Q����;�V��t��tS�d$ ������������u�[^��������̋L$U�l$;�vxS�\$V�W�D$��I �t$;���w$��    �L$$WVQ�T$,����~���;�v�L$;����t&��t"��+͋�����������u�\$�L$+�;�w�_^[]���������́�   S��$  ��W��$  uD��t@�4?  _�    [��   �D$    �D$    �D$    �D$    �D$    騽��V��$  ��wA��>  ^_�    [��   �D$    �D$    �D$    �D$    �D$    �[�����$   uA�>  ^_�    [��   �D$    �D$    �D$    �D$    �D$    �������j  �������D$    �\$�|$U��+�3�������w ��$$  ��$   PQVWS�0�������  ��$$  ����Ë�VSU��$,  ����~��$  �΋������WSU��$,  ����~��$  �ϋ�����WVU��$,  ����~��$  �ϋ�������I ;�v,�$  ;�s!VSU��$,  ����~�;�w,�
��$    �I �$  ;\$wVSU��$,  ����~��+�$  ;�vVWU��$,  �����;�wE��$  ��t+��+��(�T$��(�T$�������uዬ$$  ;��R������K����$  ;�s +�$  ;�vVWU��$,  ����t�;�r +�$  �D$;�vVWU��$,  ����t��D$�T$�ʋ�+�+�;�|2;�s�L$�D� ����   ���L$;�sF�|$��$  �\$����;�s�L$�\� ����   ���L$;�s�\$��$  �|$�������$  �D$���D$x�T� ����   �T$�D$��������]^_[��   �������������̋L$U�l$;�vxS�\$V�W�D$��I �t$;���w��    WV�T$(����~���;�v�L$;����t+��t'��+͍�$    ����������u�\$�L$+�;�w�_^[]���������́�   S��$  ��V��$  u*��t&�$;  j j j j j �    边����^[��   �U��$  ��v
��$   u'��:  j j j j j �    肹����]^[��   Ã��  �������D$    �\$�t$W��+�3�������w=��$   PUVS�������D$���D$��  �T� ����   �T$�D$���������Ë�WS��$(  ����~�Ջϋ�����VS��$(  ����~�Ջ΋�����VW��$(  ����~�Ջ΋��������    ;�v�;�sWS��$(  ����~�;�w���;\$wWS��$(  ����~�+�;�vWV��$(  �����;�wC�͋�t.��+�d$ �(�T$��(�T$�������uዬ$  ;��r������k����;�s%��I +�;�vWV��$(  ����t�;�r ��    �D$+�;�vWV��$(  ����t�D$�T$�ʋ�+�+�;�|/;�s�L$�D� ����   ���L$;��f����t$�\$�6���;�s�L$�\� ����   ���L$;��7����\$�t$����_]^[��   ���������̃=�� ���  ���\$�D$%�  =�  u�<$f�$f��f���d$���  � �~D$f(��f(�f(�f(�f(�fs�fs�5fs�4fT%��f~�f�ЋL$f��f��f~�=�  |=2   f�	�\�fV�f�t$�D$�f�!�D$�=�  �~D$tf���   ��|���f(��X�f�fT��f���f�� fT�fVĺ�  �� uf�D$�D$Ã�fD$�T$�ԃ��T$���T$���$�}  �D$����������̃=�� ��  ���\$�D$%�  =�  u�<$f�$f��f���d$�N�  � �~D$f(�f(�f(�fs�4f~�fT0�f��f�ʩ   tL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�|  ���D$��~D$f��f(�f��=�  |%=2  �fT ��X�f�L$�D$��@��f� �fT �f�\$�D$���̺j3�G�  ��3����3��j3�\�  ��3����3��=�� ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�	�  ��=�� t2���\$�D$%�  =�  u�<$f�$f��f���d$u��  ���$�24  �   ��ÍT$��3  R��<$tL�D$f�<$t�-H��  �t^�   �uA������=P� ��3  � !�   ��3  �   �u�ԩ�� u�|$ u%   �t����-�&�   �"�H3  ���� uŃ|$ u����-*)�   �=P� ��3  � !�   �2  ZËL$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+��Pd�5    �D$+d$SVW�(��  3�P�u��E������E�d�    �Pd�5    �D$+d$SVW�(��  3�P�e��u��E������E�d�    ��9  �t$�f7  �50!�  h�   �Ѓ��hX��h ��thH�P�d ��t�t$����t$�����Y�t$�l �j��_  Y�j��^  Y�V������t�Ѓ�;t$r�^�V�t$3����u���t�у�;t$r�^ËL$V3�;�u��2  VVVVV�    虱����jX^áx�;�tډ3�^ËD$V3�;�u��2  VVVVV�    �b�����jX^�95x�tۋ���3�^Ã=8� th8����  ��Yt�t$�8�Y��-  hd#hL#�6�����YYuTVWh7�\����h!�ƿH#;�Ys���t�Ѓ�;�r�=�� _^th���b�  ��Ytj jj ���3��jhH��vZ  j�k^  Y3��}�3�C9��t~����E���9}u[�5����  �E��5����  YY���u�9}�t&���u�;u�r�> t��>�  ;�t�W�  Y����ht#�h#�2���Yh|#�x#�"���Y�E������   �} u(���j��\  Y�u�����3�C�} tj��\  Y���Y  �j j�t$�������jj j �������V�  ��V�h  V��  V蒮��V�}6  V���  V���  V��W  V�  hD��h  ��$�0!^�U����u�M������E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap���jj �t$�t$�������jj �t$j �������j�]  ��Yu���ËL$�` �=�� �t�Ȟ�A�����Ȟ3�Ã|$ tZ�=�� uhD  �  ��Y���u3�áĞ��tP�H!�%Ğ �5���t$�L ����Ğt̡����,��5���5Ğ�p ��u��5Ğ�H!�%Ğ �U����e� �e� S�؅�u�����  V�u��<\t</t<:tK;�vCSV��  YY��;�u݀;:u�F;�tV�����Y�  �<\t</t<:u��+�@�E�WV�������Y�E��T  �=Ȟ�}�hh��u���  ��YY��   hd��u��n�  ��YY��   �<\t/<:t+</t'�u����  ��Y�EtP�W�����Y��   �����   �u������Y�M��ɍt|���s�;�r�jV��  ����YYt��u��uVW�n�  ����t3�PPPPP�������E��u�+��VP�l  ����t3�PPPPP�ë����W�������Y�r����}��E�uj �������Y�E������9E�tA��t�w��5����t*�!�6�7���  ��YY}�������u�v�~��u�3��V�X���Y_^[��V�5��W3��=Ȟ�=���+��hl�P��  ;�YY�6t������������Yu��9>uѡ��3��	����^�@F;�u��FPj�   ;�YYt�5���5��;������t���I��;�u�;��8��t�vP����;�Y��u��5��3�_^�VW3��t$�<�������Yu'9̞vV�t ���  ;̞v��������uɋ�_^�VW3�j �t$�t$�
���������u'9̞vV�t ���  ;̞v��������u���_^�VW3��t$�t$�!�������YYu-9D$t'9̞vV�t ���  ;̞v��������u���_^�-�  t"��t��tHt3�ø  ø  ø  ø  �SUVW�  ��U3��^WS������~�~�~3��~����8!��+Ɗ�CMu���  �   ��ANu�_^][�U��$d�����  �  3ŉ��  SW�E�P�v�x ���   ��   3����  @;�r�E���ƅ�   t+�]����;�w+�@P���  j R�I�����C�C��u�j �v�E��vPW���  Pjj ��  3�S�v���  WPW���  PW�vS�g�  ��DS�v���  WPW���  Ph   �vS�B�  ��$3��LE���t�L���  ���t�L ���  ��  �Ƅ   @;�r��M��  �E�����3�)E��U���  ЍZ ��w�L�р� ���w�L �р� ���  A;�rŋ��  _3�[蔤���Ŝ  ��jhh��jR  �"  ����,�Gpt�l t�wh��uj ����Y���R  �j�1V  Y�e� �wh�u�;5`%t6��tV�� ��u��8!tV躹��Y�`%�Gh�5`%�u�V�| �E������   뎋u�j��T  Y�U���S3�S�M���������Оu�О   �� 8]�tE�M��ap��<���u�О   �� �ۃ��u�E��@�О   ��8]�t�E��`p���[��U��� �  3ŉE�S�]V�uW�h�����3�;��}u�������3��  �u�3�9�h%��   �E��0=�   r����  �f  ����  �Z  ��P�� ���H  �E�PW�x ���)  h  �CVP�s���3�B��9U�{�s��   �}� ��   �u�����   �F����   h  �CVP�,����M��k�0�u���x%�u��*�F��t(�>����E���d%D;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   ����j�C�C��l%Zf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�.����C�S��s3��{����95О�b�������M�_^3�[藡����jh���sO  �M���'  ���}�������_h�u�����E;C�W  h   �����Y�؅��F  ��   �wh���# S�u�����YY�E�����   �u��vh�� ��u�Fh=8!tP褶��Y�^hS�=| ���Fp��   ��,��   j��R  Y�e� �C����C���C��3��E��}f�LCf�EԞ@��3��E�=  }�L��X#@��3��E�=   }��  ��`$@���5`%�� ��u�`%=8!tP����Y�`%S���E������   �0j�;Q  Y��%���u ��8!tS赵��Y�}%  �    ��e� �E��+N  Ã=�� uj��V���Y���   3��jh���M  j�Q  Y�e� �u�N��t/�����E��t9u,�H�JP�9���Y�v�0���Y�f �E������
   �M  Ë���j�}P  Y���̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t�����x�靟��V���x�菟���D$tV�"e��Y��^� VW�|$�G��tI�P�: tA�t$�N;�t��QR�!�����YYt3��%�t�t�D$� �t�t�t�t�3�@_^ËD$� � =MOC�t=csm�u+��  ���    ��  ��  ���    ~��  �   �3��jh����K  �}�]��   �s��s�u��  �   � �e� ;ute���~;w|��  �����Oȋ1�u��E�   �y t�sh  S�O�t��  �e� ��u��2���YËe�e� �}�]�u��u���E������   ;ut�w  �s�K  Ë]�u���  ���    ~��  �   �Ë �8csm�u8�xu2�H�� �t��!�t��"�u�x u�  3�A��  ���3��jh����J  �M��t*�9csm�u"�A��t�@��t�e� P�q�"����E�������J  �3�8E��Ëe��h  �L$�V�t$ƃy |�Q�I�42���^�U�����u
�  �/  �e� �? �E� ~SSV�E�@�@��ۍp~3�E����E�M�q�P�GE�P�n�������u
K�������E��E��E�;|�^[�E���j�l��u����  ���    t��  �e� ��  �M���  �n  �Mj j ���   �����j,hh��I  �ً}�u�]�e� �G��E��v�E�P蔚��YY�E��$  ���   �E��  ���   �E��  ���   ��  �M���   �e� 3�@�E�E��u�uS�uW�Қ�����E�e� �o�E������Ëe��  ��   �u�}�~�   �O��O�^�e� �E�;Fsk�ËP;�~@;H;�F�L�QVj W�������e� �e� �u�E������E    �   �E���H  ��E�맋}�u�E܉G��u��֙��Y�!  �Mԉ��   �  �MЉ��   �>csm�uB�~u<�F= �t=!�t="�u$�}� u�}� t�v�^���Y��t�uV�,���YY�jh����G  3҉U�E�H;��X  8Q�O  �H;�u�    ��<  � �u��x�t1�U�3�CS�tA�}�w��  YY����   SV�v�  YY����   �G��M��QP�����YY���   �}�E�p�tH�?�  YY����   SV�.�  YY����   �w�E�pV�n��������   ���t|��W�9Wu8���  YY��taSV���  YY��tT�w��W�E�p�e���YYPV�������9��  YY��t)SV��  YY��t�w��  Y��t�j X��@�E����  �E������E��3�@Ëe��n  3���F  �jh���wF  �E�    �t�]�
�H�U�\�e� �uVP�u�}W�F�����HtHu4j�FP�w����YYP�vS褔����FP�w����YYP�vS芔���E������DF  �3�@Ëe���  U��} t�uSV�u�Y������}  �uuV��u �K����7�u�uV�����Gh   �u@�u�F�u�KV�u�������(��tVP�ד��]�U��QQV�u�>  ���   W�(  ���    t?�  ���   ��  9t+�>MOC�t#�u$�u �u�u�u�uV�l���������   �}� u�D  �u�E�P�E�PV�u W谕�����E���;E�s[S;7|G;wB�G�O����H��t�y u*�X��@u"�u$�u�u j �u�u�u�u�����u���E��E���;E�r�[_^��U���,�MS�]�C=�   VW�E� �I��I����M�|;�|�
  �u�csm�9>��  �~� ��)  �F;�t=!�t="��  �~ �  ��  ���    ��  ��  ���   �u�  ���   jV�E���  ��YYu�	
  9>u&�~u �F;�t=!�t="�u�~ u��	  �h  ���    ��   �V  ���   �K  �u3����   ������Yu\3�9~�G�Lhd&薑����uF��;7|��4	  j�u�n���YY�EP�M��E���h���h���E�P�E�x�胙���u�csm�9>��  �~�~  �F;�t=!�t="��e  �}� ��   �E�P�E�P�u��u W�y��������E�;E���   �E�9��   ;G|�G�E�G���E�~l�F�@�X� ���E�~#�v�P�u�E����������u�M��9E���M�E��}� ��(�u$�]��u �E��u��u�u�uV�u�@����u���E����]����}�} t
jV�7���YY�}� ��   �%���=!���   �����   V������Y��   �  �  �  ���   �{  �}$ �M���   Vu�u��u$�'����uj�V�u�u�������v�����]�{ v&�} �����u$�u �u�S�u�u�uV������� �  ���    t�r  _^[��V�t$��趓���x���^� U��SVW��  ��   �E�M�csm�����"�u �;�t��&  �t�#�;�r
�@ ��   �Aft#�x ��   �} u}j�P�u�u�������j�x u�#ց�!�rX�x tR99u2�yr,9Yv'�Q�R��t�u$V�u �uP�u�u�uQ�҃� ��u �u�u$P�u�u�uQ������ 3�@_^[]�U��QQSV3��E�F3�P�u��]�������}�Y~���BWS�h �p<�f9^�F�|0v#Wh��������YYt�FC��(;�r���e� �E�_^[��V�5�&�5� �օ�t!��&���tP�5�&���Ѕ�t���  �&h���h ����t#�J�����th��V�d ��t
�t$�ЉD$�D$^�j ����Y�V�5�&�5� �օ�t!��&���tP�5�&���Ѕ�t���  �&h���h ����t#�������th��V�d ��t
�t$�ЉD$�D$^��� � V�5�&�� ����u�5���k���Y��V�5�&�� ��^á�&���tP�5 ��A���Y�Ѓ�&���&���tP�� ��&��HA  jh��m>  h���h �E�u�F\�)3�G�~��t/������t&h���u�d �Ӊ��  h���u��Ӊ��  �~pƆ�   CƆK  C�8!�FhP�| j��A  Y�e� �E�Fl��u��-�Fl�vl�v  Y�E������   �	>  �j��@  Y�VW�D �5�&�������Ћ���uNh  j�z�������YYt:V�5�&�5������Y�Ѕ�tj V�����YY�, �N���	V����Y3�W�� _��^�V��������uj� ���Y��^�jh(��=  �u����   �F$��tP輤��Y�F,��tP认��Y�F4��tP蠤��Y�F<��tP蒤��Y�FD��tP脤��Y�FH��tP�v���Y�F\=�)tP�e���Yj�@  Y�e� �~h��tW�� ��u��8!tW�8���Y�E������W   j�k@  Y�E�   �~l��t#W�u  Y;=�-t���,t�? uW�s  Y�E������   V����Y�j<  � �uj�<?  YËuj�0?  YÃ=�&�tLW�|$��u&V�5�&�5� �օ�t�5�&�5�&���Ћ�^j �5�&�5���`���Y��W����_��&���t	j P�� �Wh���h ����u	�����3�_�V�5d h��W��h��W�����h��W�����h��W����փ=�� �5� � �t�=�� t�=�� t��u$�� ����� ������5��� ��� �����&��   �5��P�օ���   �X����5��������5�����������5�����������5 ������������ ��=  ��teh���5������Y�Ѓ����&tHh  j�L�������YYt4V�5�&�5�������Y�Ѕ�tj V�����YY�, �N��3�@��l���3�^_�jhP��:  ������@x��t�e� ���3�@Ëe��E������  �*:  ������@|��t������jhp���9  �5��[���Y��t�e� ���3�@Ëe��E������}���h������Y��������U���SQ�E���E��EU�u�M�m��]�  VW��_^��]�MU���   u�   Q�;�  ]Y[�� U���(  ���������5 ��=��f�(�f��f���f���f�%�f�-��� ��E ���E���E�$��������`�  ������	 ���   �  �������$ �������$ �X�j�4  Yj �  h��� �=X� uj�  Yh	 �� P� �ËL$S3�;�VWt�|$;�w�  j^�0SSSSS�=��������1�t$;�u��ًъ�BF:�tOu�;�u��a  j"Y�����3�_^[�U���V�u�M�蟬���u�P�Y�����e�F�P�J�  ��Yu��P�<�����xYuFF�M����   �	��	�F�����F��u�8M�^t�E��`p���U���V�u�M��.����E��ɋu�t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B�Ɉu��}� ^t�E��`p�����D$�����Az3�@�3��U��QQ�} �u�ut�E�P��  �M��E��M��H��EP��  �E�M�����j �t$�t$�t$������Å�V��tV�@���@PV�V蕍����^�j �t$�z���YY�j �t$�����YY�U���SVW�u�M�������3�;�u+�  j_VVVVV�8�:������}� t�E��`p����!  9uv�9u~�E�3���	9Ew	�V  j"뺀} t�U3�9u��3Ƀ:-����ˋ��:����}�?-��u�-�s�} ~�F�����E����   � � �3�8E��E��}�u����+�]h��SV� �����3ۅ�tSSSSS�w�����9]�Nt�E�GF�80t.�GHy���-F��d|
�jd_�� ��F��
|
�j
_�� �� F�L�t�90uj�APQ�������}� t�E��`p�3�_^[��U���,�  3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�1�  3ۃ�;�u�  SSSSS�0贊�������o�E;�v����uu����3Ƀ}�-��+�3�;���+��M�Q�NQP3��}�-��3�;�����Q�M�  ��;�t���u�E�SP�u��V�u��������M�_^3�[������U��j �u�u�u�u�u������]�U���$VW�u�M��E��  3��E�0   螨��9}}�}�u;�u+�+  j^WWWWW�0�ˉ�����}� t�E�`p����  9}vЋE��9E� w	��
  j"���}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW� �������t�}� � ��  �M�ap��  �;-u�-F�0F�} je����$�x�FV��  ��YY�L  �} ���ɀ����p��@ �2  %   �3��t�-F�]�0F������$�x��OF��ۃ����  �3���'3��u!�0�O����� F�u�U���E��  ��1F��F9U�Eu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~M�W#U���M�#E���� ���  f0 ��f=9 vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� ��  f= v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V������u�E�8 u���} �4����$�p���WF�4�  3�%�  #�+E�SY�x;�r�+F�
�-F�����;Ӌ��0|$��  ;�rSQRP��  0�F;��U�����u��|��drj jdRP���  0��U�F����;�u��|��
rj j
RP���  0��U�F���]�0��F �}� t�E�`p�3�[_^��U���SVW�u�؋s���M�N�4�����u-��  j^�03�PPPPP�j������}� t�E��`p����   �} v̀} t;uu3��;-����� 0�@ �;-��u�-�w�C3�G�����n����0F���} ~D���Y����E����   � � ��[F��}&�ۀ} u9]|�]�}���(���Wj0V�L������}� t�E��`p�3�_^[��U���,�  3ŉE��ESVW�}j^V�M�Q�M�Q�p�0���  3ۃ�;�u�  SSSSS�0�b��������Z�E;�v���u��3Ƀ}�-��+��u�M�Q�M��QP3��}�-���P��  ��;�t���u�E�SV�u���d������M�_^3�[�؀����U���0�  3ŉE��ESV�uWj_W�M�Q�M�Q�p�0�&�  3ۃ�;�u�  SSSSS�8詄�������   �M;�vދE�H�E�3��}�-������<0u��+ȍE�P�uQW�W�  ��;�t��X�E�H9E������|-;E}(:�t
�G��u��_��u�E�j�u���u��������u�E�jP�u���u�u�������M�_^3�[������U��E��et_��EtZ��fu�u �u�u�u�u�&�����]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u������u �u�u�u�u�u�|�����]�U��j �u�u�u�u�u�u�^�����]�VW3����&�6�:�������(Y�r�_^�Vh   h   3�V�#�  ����tVVVVV������^�U������]����]��E��u��M��m��]����]�����z3�@��3���h4��h ��th�P�d ��tj ��������zuf��\���������?�f�?f��^���٭^�����&�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�����&�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp�����&���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-�&��p��� ƅp���
��
�t���������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR��  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   ��@��   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z��l������������\������   s��|���d������������T������   v��t�떋D$3�;��&tA��-r�H��wjXË��&�D���jY;��#����������u�X(Ã��������u�\(Ã��V������L$Q�����Y��������0^Ã%�� �U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]Ã%�� �)�  ���3��U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]�U��$X�����(  �  3ŉ��  �`(Vtj
��   Y�o�  ��tj�q�  Y�`(��   ���   ���   ���   �]|�ux�}tf���   f���   f�]pf�Elf�ehf�md����   ���  ���  ���   �E�  ���   �@�jP���   �E�j P��{���E����EЍE�j �E�  @�u��E��  �E�P� j�;���̋L$�`(�T$#T$��#�ʉ`(�QS�\$VW3�3�;�h(tG��r���w  Uj�Ⱦ  ��Y�1  j跾  ��Yu�=l��  ���   �?  h(��  S�0�U��������tVVVVV�py����h  �I�Vj �M� �� ��u&h�h�  V���������t3�PPPPP�,y����V�����@��<Yv8V������;�j�D�h�+�QP�K�  ����t3�VVVVV��x�����3�h�SU贼  ����tVVVVV��x�����4�l(SU蒼  ����tVVVVV�x����h  h��U豺  ���3j��� ��;�t%���t j �D$P�4�l(�6�	���YP�6U�� ]_^[Y�j�M�  ��Ytj�@�  ��Yu�=l�uh�   �4���h�   �*���YYËD$�L�������U���������$�\$�   ��fD$f=�f�fT���fs�,f�� fV�f��%�   ��%�  �Y<�P�f,�P��f(4�`���  +у�ʁ�   ���  �    �� fn�f��fs����f8��fs�&f�� fT%�%�   ��%�  �Y�p��Y,�p��fX4���fV%��X�fT���fs�f�� f8�\�f=@%�  ��%�  �Y,����Y���fX4ŠfT��\��X����Y��Y��Y��\��Y����\��X�fL$f���\��\�f8f���\����X��\��\�f�%�  =�  �  ���  -�?  º�@  +�-p<  Ё�   ���  �\��\�f%8fT�fT��\�fWҺ`@  f�����Y��\��\��Y��Y�f(��Y��-��Y�f(��X�fp���X�� +��� �-�� �� ��  ȃ��ခ��� �X����X�fY��\�fY��\�����f(��f(5fY�fX�fp���Y�fW���?  �X�f���X�f%0fn��YT$�Y�fs�-fp�Df(= �X�fY��X�f�fY��Y�fY�fX�fY��Y�fp���Y�fp���Y��Y��XŃ��X��X��X�fD$�D$���fL$f f~���fT�fs� f~Ɂ�  ���   ��� �  �� �  �ځ��  fs�4fVӹ�  fn�fs�f��f��f��f��fv�f�ʁ��  ���  ��  %�   =�   ��  fL$fT$��  fn�fT fs�4f��f`f��fv�f��%�   �� ȁ�   ��r^�� f�f��&���f|$fd$f~�fs� f~���%���=  ���  ��  �� ��  �  �    fW���C  f��f=�f��Y�f~�fs� f~��� tRfT���fT fs�,f�� fV�%�   ��%�  �Y<�P�f,�P��f(4�`��> �\����Ё������ u��T$��   ��� t1��#��  ��fn�fs� f�fT$�^ʺ   �  ��#��� ��   ���f�fW�fT�fv�f�Ɂ��   ���   ��   f���� �  �� ��   %�   =�   uefL$fT$��  fn�fT fs�4f��f��f��fv�f��%�   =�   t#fL$f��% �  �� t�`��X�fL$f��% �  �� �G  ���fL$f��% �  �� �+  ����X��ĺ�  �  fT$f~�fs� f~ҁ����¹    �� �����fHf��Yɺ   �H  fd$fT$f�fW�fT�fv�f��%�   =�   ��   f~��� u fs� f~��  �?��   ��  �u���f�fW�fT�fv�f��%�   =�   uUf��fd$% �  ��  �у� ��   �� tf��%�  =�?  r���f��%�  =�?  s����P��X��º�  �cf~�fs� f~��������f��   �� t:f~�   %���=  �w%r�� w��fD$�D$���fP��   ��fD$�T$�ԃ��T$���T$���$�@8  �D$��Ã� ~(=   �<  V�Ѓ��� � ��   ��W��?  �&= ����  V�Ѓ����   � � W�    �X����X����� fY��\�fY��\�����f(��f(5fY�fX�fp���Y��X��X�f%0fnʁ�� �������� �fW���?  f���YT$�Y�fs�-fp�Df(= �X�fY��X�f�fY��Y�fY�fX�fY��Y�fp���Y�fp���Y��Y�fn�fs�-fn�fv�f���X��X�fT��X�fW�fv�f���\����X�fT�f��_�\��X��XÃ� N^�Y��Y��X��Y��X�f��%�  �   =�  �����   �� ������fD$�D$���^�X��Y��Y��X�f��%�  �   =�  ������   �� �������fD$�D$���fxfn��Y�fs�-fV��   �����   �� tfh�Yp�e���fp�Y��T���fp�DfY�f��%�  ��@  +�-p<  Ё�   ������=   �r �ɀ� fn�fs�-��fD$�D$���fd$f�����  ���?  f��3�% �  �� �-����K�����$    ��$    �ƅp����
�uK�����ƅp����2������;  ������a���t��=T�t����=H  ��@u��
�t�������F  �t2��t������������.��������- )ƅp����������ݽ`������a���Au����ƅp������-*)�
�uS��������
�u�����>�����   ����
�u���u
�t���ƅp����- )��u�
�t������������������X��ݽ`������a���u���- )
�t���ƅp�������������- )ƅp����
�u����- )������->)�ٛݽ`������a���Au�������ݽ`������a���������ݽ`�������������ٛ���u���R)�����ٛ���t�   ø    ���   ��V��t��V���$���$��v�z   ���f���t^��t�����U��QQ�EQQ�$��  ��YYuH�EQQ�$�Ư  �]YY����Dz/�EQ��$Q�]��E��$衯  �]�YY����DzjX��3�@��3���U����V�U3�3����E��Au��  �9E�  ��u=9Uu��������z�������(2��   ��������A�Eu����   ����   9MuB9Uu=��������z	�����   ���������Ez�(2�   �023��F�   9E��u&9Uu�U�����v����U����A�EtZ�����T9M��uY9UuT�EQQ�$������Y�UY������z�����(2u����U����Au��u���H2�E���������؋�^]�U��QV�uV�!����E�F��Yu�0���� 	   �N ����-  �@t����� "   ��S3ۨt��^��   �N�����F�F����f��F�^�]�u,�
_  �� ;�t��^  ��@;�u�u�®  ��YuV�s�  Yf�FW��   �F�>�H��N+�I;��N~WP�u�=x  ���E��M�� �F����y�M���t���t����k�8����������)�@ tjSSQ�q  #����t%�F�M��3�GW�EP�u��w  ���E�9}�t	�N �����E%�   _[^��U��$�����x  �  3ŉ��  ��   S��  V3�W��  ��  �M��EЉ}ԉu��u�u��u��uĉu��u�����9u�u-����VVVV�    V�(h�����}� t�E��`p������  �E��@@��   P�/������Yt6�u��!������Yt(�u������u����4���������k�8YY3����)�@$�u����u��܆�����Yt6�u��Ά�����Yt(�u�������u����4���讆����k�8YY3����)�@$��"���;������3Ʉ҉ủu؉u��U���  C�}� �]���  ��, <Xw�������3��3�3�����j��Y;��E��z  �$��0�M���u��u��u��uĉu�u��X  �� t>��t-��tHHt���9  �M��0  �M��'  �M��  �M�   �  �M��	  ��*u ���}ԋ�;��}���  �M��]���  �E�k�
�ʍDЉE���  �u���  ��*u���}ԋ�;��}���  �M���  �E�k�
�ʍDЉE��  ��ItF��ht8��lt��w�x  �M�   �l  �;luC�M�   �]��W  �M��N  �M� �E  �<6u�{4uCC�M� �  �]��(  <3u�{2uCC�e�����]��  <d�  <i��  <o��  <u��  <x��  <X��  �u��E�P��P�u��~M  Y���E�Yt�MЍu���  �C���]���  �MЍu���  �  ��d�r  ��  ��S��   tZ��AtHHt@HHtHH�N  �� �E�   �U�M�@9u��]�   �]܉E���  �E�   �	  f�E�0uu�M�   �lf�E�0u�M�   �M����u������f�E��}ԋ��}���  ;�u��)�E܋E��E�   �  ��X�9  HHt]+��d���HH��  ��f�E��}�t'�G�Ph   �E�P�E�P�)�  ����t�E�   ��G��E��E�   �E�E��P  ���;Ɖ}�t.�H;�t'f�E� � �M�t�+����E�   �  �u��  �|)�E�P�K���Y��  ��p��  �t  ��e��  ��g�������itY��nt��o��  �E��E�   tI�M�   �@�7���}�舠������  �E� t	f�E�f���Ẻ�E�   �  �M�@�E�
   �M�f���C  ��W���k  u��guG�E�   �>9E�~�E��}�   ~-�u���]  V�?������U�Y�E�t
�E܉u�����E�   3�����E��G��E��E�P�u����u��}�P�u��E�SP�5�&�����Y�Ћ}����   t9u�u�E�PS�5�&�����Y��YY�}�gu;�u�E�PS�5�&����Y��YY�;-u�M�   C�]�S�r����E�   �M��!��s�p���HH��������Y  �E�'   �E��E�   ������E�Q�E�0�E��E�   ����f�� ��������� t��@�}�t�G���G�����@�G�t��3҉}���@t;�|;�s�؃� �ځM�   f�E� ��ڋ�u3ۃ}� }	�E�   ��e���   9E�~�E����u!Eč��  �E��M������t$�EؙRPSW�M�  ��0��9�]�����~M��N�̍��  +�Ff�E� �E؉u�tL��t�΀90tA�M܋M��0@�2If90t@@;�u�+E����;�u�|)�E܋E��I�8 t@;�u�+E܉E؃}� ��   �E�@t%f� t�E�-��t�E�+��t�E� �E�   �]�+]�+]��E�u�uЍE�Sj �H�  ���uċ}ЍE̍M��X�  �E�Yt�E�uWSj0�E���  ���}� �E�tQ��~M�u܉E���M�Pj���  P�E�FPF� �  ����u9E�t�u��E̍��  ��  �}� Yu���M����M�P�E��֧  Y�}� |�E�tWSj �E�虧  ���}� t�u��	q���e� Y�]�����E�t$�M��}Ԋ��)��������    3�PPPPP�$����}� t�E��`p��E̋��  _^3�[�[�����  �û*")=)�)�)�)*�*U��� S3�9]u �G���SSSSS�    ��^��������   V�uW�};�t!;�u����SSSSS�    �^��������j����;��E�w�}��u�E��u�E�B   �u�u�P�u��U��;�Et4;�|"�M�x�E����E�PS�a������YYt�E�3�9]�\>���HH_^[��U��S3�9]u����SSSSS�    �^��������[V�u;�t9]w�V����    �0�u�u�u�uVh���������;�}����u�$���� "   SSSSS��]�������^[]�jTh���{  3��}��E�P�L!�E�����j8j ^V�C���YY;��   ����5d���   �)�@ ���@
�x�@$ �@%
�@&
��8�����   ;�r�f9}���   �E�;���   �8�X�;�E�   ;�|��3�F�Rj8j �����YY��tM������d� ��   �&�@ ���@
�` �`$��@%
�@&
��8���   ;�r�F9=d�|���=d��e� ��~m�E����tV���tQ��tK�uQ�H ��t<�u�������k�84����E� ���Fh�  �FP�؍  YY����   �F�E�C�E�9}�|�3ۋ�k�85������t���t�N��r�F���uj�X�
��H������P�� �����tC��t?W�H ��t4�>%�   ��u�N@�	��u�Nh�  �FP�B�  YY��t7�F�
�N@�����C���g����5d��� 3��3�@Ëe��E���������  �VW����>��t1��   �� t
�GP�\ ���8   ;�r��6��l���& Y������|�_^�S3�9��VWu�����5`�3�;�u����   <=tGV覧��Y�t�:�u�jGW蟯����;�YY�=��tˋ5`�U�@V�u�����E�>=Yt/jU�q���;�YY�tJVUP�D�������tSSSSS�Y�������8u��5`��l���`�����   3�Y]_^[��5����k����������QQ�P�SUVW�=� 3�3�;�j]u-�׋�;�t�P�   �"�D ��xu	�ţP���P�����   ;�u�׋�;�u3���   f9��t�f9u��f9u�=� SSS+�S��@PVSS�D$4�׋�;�t2U�*���;�Y�D$t#SSUP�t$$VSS�ׅ�u�t$�k��Y�\$�\$V�� ���X;�t;�u��� ��;��p���8t
@8u�@8u�+�@��U�­����;�YuV�� �D���UVW��]����V�� ��_^][YY�VW����;ǋ�s���t�Ѓ�;�r�_^�VW����;ǋ�s���t�Ѓ�;�r�_^�U��QQV�E�3�P�u��u�������YtVVVVV�W�����E�P�!�����YtVVVVV�W�����}�^u�}�r3�@��jX��3�9D$j ��h   P�� ���T�u3���}������`�u$h�  �9  ��Yu�5T��� �%T� ��3�@�U3�=`�uTS�4 W3�9-H�~1V�5L���h �  U�v��� �6U�5T��Ӄ�G;=H�|�^�5L�U�5T���_[�5T��� �-T�]��U��QQV���������F  �V\�L*W�}��S99t��k����;�r�k��;�s99u���3���t
�X�ۉ]�u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   �@*�=D*���;�}$k��~\�d9 �=@*�D*B߃�;�|�]�� =�  ��~du	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�øcsm�9D$u�t$P����YY�3��h@:d�5    �D$�l$�l$+�SVW�  1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q���̃�S�\$ UV�s35  W�����D$ �D$   �{t�N�38�Q���N�F�38�rQ���D$(�@f�  �k����L$0�T$�D$�L$ �S�t^�Dm �L��ɍ\���D$t���hX  ���D$|DL�D$�����ù|$ t$����t�N�38��P���N�F�38��P���D$_^][����D$    �ƋL$(�9csm�u*�=p� t!hp��l�  ����t�T$(jR�p����L$,�X  �D$,9hth  W�Ջ��X  �D$,�L$�H����t�N�38�_P���N�V�3:�OP���K���W  �{��P���h  W�˺�����W  ����U����  �e� �e� SW�N�@�;ǻ  ��t��t	�У$ �`V�E�P�` �u�3u��� 3��, 3��� 3��E�P�� �E�3E�3�;�u�O�@����u������5  �։5$ ^_[��VW3��X��<�T*u��P*�8h�  �0����  ��YYtF��$|�3�@_^Ã$�P* 3���S�\ V�P*W�>��t�~tW��W��d���& Y����p+|ܾP*_���t	�~uP�Ӄ���p+|�^[�U��E�4�P*�� ]�jh������3�G�}�3�9T�u����j�����h�   诠��YY�u�4�P*9t���nj�#���Y��;�u������    3��Qj
�Y   Y�]�9u,h�  W���  YY��uW��c��Y�����    �]���>�W��c��Y�E������	   �E��S����j
�*���Y�U��EV�4�P*�> uP�$�����Yuj诟��Y�6�� ^]�h@  j �5T��< ���L�uËL$�%�� �%H� �T�3��P��X�   @ËH��L�k����T$+P��   r	��;�r�3��U����M�AV�uW��+y�������i�  ��D  �M��I���M���  S�1��U�V��U��U����]ut��J��?vj?Z�K;KuB�� �   �s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J;։M�v��;�t^�M�q;qu;�� �   �s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���� �Ls%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   �������   �\��5� h @  ��H� �  SQ�֋\�����   ���	P����@�\�����    ����@�HC����H�yC u	�`�����x�ueSj �p�֡���pj �5T��4 �H����k��L�+ȍL�Q�HQP�O���E���H�;��v�m�L��T��E����=\�[_^�áX�V�5H�W3�;�u4��k�P�5L�W�5T��P ;�u3��x�X��5H��L�k�5L�h�A  j�5T��< ;ǉFt�jh    h   W�� ;ǉFu�vW�5T��4 뛃N��>�~�H��F����_^�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W�� ��u����   �� p  ;��U�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[��U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I��?�M�vj?Y�M��_;_uC�� �   �s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O��?�L1�vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���� �Ls�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N��?�]�K�vj?^�E���   �u���N��?vj?^�O;OuB�� �   �s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���� �Ls�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[��U����H��Mk�L�������M���SI�� VW}�����M���������3���U��T�����S�;#U�#��u
��;؉]r�;�u�L���S�;#U�#��u
��;ى]r�;�u[��{ u
���];�r�;�u1�L��	�{ u
��;ى]r�;�u�����؅ۉ]u3��	  S�@���Y�K��C�8�t�T��C�����U�t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��ɍy�>u;��u�M�;\�u�%�� �M���B_^[�ËD$�����5���`�����Yt�t$�Ѕ�Yt3�@�3������U�������$�~$�   ��fD$f%�2f�2fW�f�2��fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU *fV�f($� ���X��\��Y��Y��Y����X��^�f=h2f-X2�\�fs�?��fs�?�Y�fp�Df5`2�Y��Y���fW��Y��Y��X��Y��X�fp���X��X��X�fD$�D$���-�  ��C�  �Y��\��Q�f��fs�fT=P2fs���f%�2���\��Y��X��\��Y���fT�fs�f��fVՁ���  ��Y<� *�Y�f( 2�Y��Y��\��X��\��X�f-X2�\��X�fh2�^�f`2f\� ���Y�%�   ���Y��Y΃��Y��Y��X�f���Y��X�f���X�fp���\��X�fV�fD$�D$����;  = 8  sjf�f(5p2f�f(�2f(%�2fY���fY�fY�fY����Y�fX�fY��Y�fX�fY�fp���X��X�fD$�D$���-�;  ���O  �Y��\��Q�f��fT=@2fp�DfT@2��f%�2���\��Y��X��Y��\����Y��Y��\��\��X��\�f(p2fp���\��X�fp���X��Y��X�fp���^�f(�2f(-�2f(�2fY���fY�fY�% �  �Y�fY�fX�f(��Y�fY�f( 2�Y�fX�fp���Y��fY��X�fW�fp���Y�fp���X���f���\��X��X��X��\��\��\��\�fV�fD$�D$����� = � ��   f~�fs� f~�����  �?+���� ��   fT$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��=   ��fD$�T$�ԃ��T$���T$�$�	  fD$����fD$�D$���f�2f 2f(2�X�fU�fV���fD$�D$���fD$fW��Xƺ�  �t���fD$fW�����f�����  �����  r�X�fV��Y�fD$�D$���U�������$�~$�   ��fD$f%�Jf�JfW�f�J��fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU BfV�f($� 3���X��\��Y��Y��Y����X��^�fxJf-hJ�\�fs�?��fs�?�Y�fp�Df5pJ�Y��Y���fW��Y�f\% J�Y��X��Y��\�fp���X��\��\�fD$�D$���-�  ��A�-  fs�&fs�&f��fU��\����Y��X�fV��\��Y����\��Q�%�   ������fT�fs�f��fV�fn�fp� ����  ��Y<� B�Y��Y��Y��\�fTJ�X��\��X�f-hJ�\��X�fxJ�^�fpJfX� 3���Y��Y��Y΃��Y��Y��X�f���Y��X��X�% �  f����fp���X��\��X��X��X�fW�fD$�D$����;  = 8  ��   f�f(5�Jf�f(�Jf(%�JfY�f(- J��fY�fY�fY����Y�fX�fY��Y�fX�fp��fY�fp���\�fp���\��\��\��\��\��X�fD$�D$���-�;  ����   fW�fT=�Jf%�Jf(�J�Y�f(�J�\�f(�Jfp�D�Q�fY�fp�Df��fY�fX�f@JfY�����Y�fX�fp�D�Y�fTJfY�fT�fp�D�\��X��Y��\��\��Y�fp���\��^��fX�fY�fp���X�% �  f��fp���X��X��X��X�fW�fD$�D$����� = � ��   f~�fs� f~�������  �?+���� ��   fT$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��:   ��fD$�T$�ԃ��T$���T$�$�  fD$����fD$�D$���f������fn�fp� f Jf(JfT�fT��X�fD$�D$���f JfJ�X�fD$�D$���fW��Xƺ�  �J���������������U�������$�~$�   ��fD$f��f%�f-00f=��B  fPS�Y�fXS�-��X�fpS�\�f(`S�Y�fɁ�v ����?f(-@S�K���fY��\��YxS�\�fxf����\�fY�f\�f(5 S�Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-0S�Y fX5SfY����XXfY����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���+f��f%�f����f�S�\�fL$�D$����O���I ����U�������$�~$�   ��fD$f��f%�f-00f=��B  f \�Y�f\�-��X�f \�\�f(\�Y�fɁ� v ����?f(-�[��S���fY��\��Y(\�\�fxf����\�fY�f\�f(5�[�Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-�[�Y fX5�[fY����XXfY����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���I��f��f=�u�Y@\fD$�D$���f0\�Y��\��Y8\fD$�D$�����N���U���(3�9��S�]V�uW�}�E��E��E��E��E��E��E��E�t�5D�订��Y��6��M��   ;��t  �[  ����   ��   ��jY+���   J��   ����   J��   ��tqJtE��	��  �E�   �E�]��M��]�Q��]���]��Ѕ�Y��  ������ "   �  �E�]��M��]�Q��E�   �]���]���Y�j  �E�   �E�]��E�]��]���]���"  �M��E�]�r����E�]�׉M��E�]�Z����E�]놃�tNIt?It0It ��t����   �E�]��E��\��E�]����E�]�x����E�   ��������   �E�   �E��\��������������   �$�Z�E�]��E�]��E�]��E��\��E��\��E��\�y����E��\�m����E��\��E��\��E��\��M����]���]�M��]�Q�E�   �Ѕ�Yu�e���� !   �E��_^[�Ë�yY�Y�Y�Y�Y�Y1Y�YYY�Y�Y�YU��QQSV���  V�5p+�D_  �EYY�؋EQf%�f=�Q�$uU�)W  ��YY~-��~��u#�ESQQ�$j��]  ���rVS��^  �EYY�d�ES��$���\$�E�$jj�?�y  �]��EY�]�Y����DzVS�^  �E�YY�"�� u��E�S���\$�E�$jj��]  ��^[���������U�������$�~<$�   ���~|$f�f(�fT0]f/X^��  �U  f/H^snf/P^��  f(�fY�f(�fY�f(- ^fY�fX-�]fY�fX-�]fY�fX-�]�Y�f(�f���X��Y��\�f�|$�D$�f/@^��   f(�fY�f(�fY�f(-�]fY�fX-�]fY�fX-�]fY�fX-�]fY�fX-�]fY�fX-p]fY�fX-`]fY�fX-P]�Y�f(�f���X��Y��\�f�|$�D$��~�fW�f/8^sO�~0^�~-^�~��X�fs�,f��f~؍@�~,���~��\��Y��X(^�^�f���   �~��~ ^�^�f��~�ؕ�~$���f(�fY�f(�fY�f(- ^fY�fX-�]fY�fX-�]fY�fX-�]�Y�f(�f���X��Y��\��\��\�fV�f�D$�D$�f/^u�D$�f/`^s�h^�h^���$�$���D$��h^�h^�D$��~��~ ]fT�f.�z�D$���h^��@]ú�  ���T$�ԃ��T$�T$�$�������D$Ð����U�������$�~$�   ��fD$�    f(�f�fs�4f�� f(p^f(�^f(%�^f(5�^fT�fV�fX�f�� %�  f(�P_f(�`cfT�f\�fY�f\��X�fY�f(�fXƁ��  �����  ��   ���  ��*�f���
��   �    �� D�f( _f(�f(0_fY�fY�fX�f(@_�Y�f(-�^fY�f(��^fT�fX�fX�fY��Y�fX�f(�f�fY˃�f(�f��X��X��X�fD$�D$���fD$f(�^��� f�� �� wH���t^���  wlfD$f(p^f(�^fT�fV���� f�� �� t�_ú�  �Of�^�^�f _�   �4f�^�Y�������/��������  ���  s:fW��^ɺ   ��fL$�T$�ԃ��T$���T$�$�Q����D$���fT$fD$f~�fs� f~с��� ��� t���  릍d$ U���0���S�ٽ\�����=�3 t�7�����8����   [����ݕz������U���U���0���S�ٽ\����=�3 t蓬����8�����8�����Z   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���ƅq���蜬���   [�À�8�����=P� uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   ��g�����������xg����s4��g�,ǅr���   ��g�����������pg����v��gVW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P��l  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8����贪������[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[���l$�l$�D$���   5   �   t��������+ u��ËD$%�  tg=�  t`�|$�D$?  %��  �D$ �l$ �D$%�  ��t��+����+���l$�����+����+���l$��ËD$D$u��ËD$%�  u��|$�D$?  %��  �D$ �l$ �D$%�  t=�  t2�D$�s*��D$�r ��������+�|$�l$�ɛ�l$������l$��Ã�,��?�$��+����,Ã�,�����,Ã�,�����,�����,�����,�����,��|$���<$�|$ �����l$ �Ƀ�,Ã�,��<$�|$�����l$�Ƀ�,Ã�,����|$���<$�|$ �^����l$ ��,��<$�|$�J�����,��|$�<$�:����l$��,��|$�<$�&�����,��|$�����<$�|$ �������l$ �ʃ�,Ã�,��<$���|$��������l$�ʃ�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$�����Ƀ�,��|$���<$�������l$��,��|$���<$�����Ƀ�,��|$�����<$�|$ �j������l$ �˃�,Ã�,��<$���|$�K������l$�˃�,Ã�,����|$�����<$�|$ �$������l$ ��,��<$���|$�����ʃ�,��|$���<$��������l$��,��|$���<$������ʃ�,��|$�����<$�|$ ��������l$ �̃�,Ã�,��<$���|$�������l$�̃�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�h����˃�,��|$���<$�T������l$��,��|$���<$�<����˃�,��|$�����<$�|$ �"������l$ �̓�,Ã�,��<$���|$�������l$�̓�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$������̃�,��|$���<$�������l$��,��|$���<$�����̃�,��|$�����<$�|$ �~������l$ �΃�,Ã�,��<$���|$�_������l$�΃�,Ã�,����|$�����<$�|$ �8������l$ ��,��<$���|$� ����̓�,��|$���<$�������l$��,��|$���<$������̓�,��|$�����<$�|$ ��������l$ �σ�,Ã�,��<$���|$�������l$�σ�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�|����΃�,��|$���<$�h������l$��,��|$���<$�P����΃�,Ã�,�<$�|$�;�����,Ã�,�|$�<$�(�����,�P�D$%  �=  �t3��% 8  t�D$����X� �Ƀ��<$�D$�����,$�Ƀ�X� �t$X� P�D$%  �=  �t3��% 8  t�D$�k���X� �Ƀ��<$�D$�V����,$�Ƀ�X� �t$X� P��% 8  t�D$�/���X� �Ƀ��<$�D$�����,$�Ƀ�X� P��% 8  t�D$�����X� �Ƀ��<$�D$������,$�Ƀ�X� P�D$%  �=  �t3��% 8  t�D$�����X� �Ƀ��<$�D$�����,$�Ƀ�X� �|$X� P�D$%  �=  �t3��% 8  t�D$�~���X� �Ƀ��<$�D$�i����,$�Ƀ�X� �|$X� P��% 8  t�D$�B���X� �Ƀ��<$�D$�-����,$�Ƀ�X� P��% 8  t�D$����X� �Ƀ��<$�D$������,$�Ƀ�X� P��,�<$�|$������,X�P��,�|$�<$�������,X�PSQ�D$5   �   ��  �������+ �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u������+�Ƀ�u�\$0�|$(���l$�-�+�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8��+�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$3ҋD$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w����+�|$��+�<$� �|$$�D$$   �D$(�l$(����+�<$�l$$�T�����0Z�����0Z�PSQ�D$5   �   ��  �������+ �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u������+�Ƀ�u�\$0�|$(���l$�-�+�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8��+�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$�    �D$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w����+�|$��+�<$� �|$$�D$$   �D$(�l$(����+�<$�l$$�Q�����0Z�����0Z�������@��������������̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[�SUV�t$���   3�;�Wto=�4th���   ;�t^9(uZ���   ;�t9(uP��/�����   �cr  YY���   ;�t9(uP��/�����   �r  YY���   ��/�����   �/��YY���   ;�tD9(u@���   -�   P�/�����   ��   +�P�/�����   +�P�x/�����   �m/�������   �=�3t9��   uP��o  �7�F/��YYj�~P[���,t�;�t9(uP�%/��Y9o�t�G;�t9(uP�/��Y��Ku�V�/��Y_^][�SUV�t$W�=| V�׋��   ��tP�׋��   ��tP�׋��   ��tP�׋��   ��tP��j�^P]�{��,t	���tP�׃{� t
�C��tP�׃�Mu؋��   �   P��_^][�V�t$��tSUW�=� V�׋��   ��tP�׋��   ��tP�׋��   ��tP�׋��   ��tP��j�^P]�{��,t	���tP�׃{� t
�C��tP�׃�Mu؋��   �   P��_][��^Å�t7��t3V�0;�t(W�8�������YtV�R����> Yu���,tV�x���Y��^�3��jh�������袈�����,�Fpt"�~l t苈���pl��uj �i��Y��������j����Y�e� �Fl�=�-�i����E��E������   ��j����Y�u��U����  3ŉE�SV3�9ܦW��u8SS3�GWh$hh   S�<!��t�=ܦ��D ��xu
�ܦ   9]~"�M�EI8t@;�u�����E+�H;E}@�E�ܦ����  ;���  ����  9] �]�u��@�E �5� 3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w��B����;�t� ��  �P�f+��;�Yt	� ��  ���E���]�9]��=  W�u��u�uj�u �օ���   �5<!SSW�u��u�u�֋�;ˉM���   f�E t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w�6B����;�tj���  ���P�*��;�Yt	� ��  �����3�;�tA�u�VW�u��u�u�<!��t"9]SSuSS��u�u�u�VS�u �� �E�V�P��Y�u��P���E�Y�Y  9]�]�]�u��@�E9] u��@�E �u�mn  ���Y�E�u3��!  ;E ��   SS�MQ�uP�u �n  ��;ÉE�tԋ58!SS�uP�u�u��;ÉE�u3��   ~=���w8��=   w� A����;�t����  ���P�)��;�Yt	� ��  �����3�;�t��u�SW�7�����u�W�u�u��u�u��;ÉE�u3��%�u�E��uPW�u �u���m  ���u������#u�W�lO��Y��u�u�u�u�u�u�8!��9]�t	�u��)��Y�E�;�t9EtP�)��Y�ƍe�_^[�M�3�������U����u�M��6���u(�M��u$�u �u�u�u�u�u�-����� �}� t�M��ap���U����u�M��l6���E�M����   �A% �  �}� t�M��ap���j �t$����YY�U���S�u�M��'6���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�u�����YYt�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�rO  �� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�ËD$��VW|Z;d�sR����k�8�����<�����<�u6�=l�S�\$u�� tHtHuSj��Sj��Sj��� ��3�[�軗��� 	   �×���  ���_^ËL$S3�;�VW|[;d�sS���k�8�����<������@t5�8�t0�=l�u+�tItIuSj��Sj��Sj��� ���3���:���� 	   �B�������_^[ËD$���u�+����  ����� 	   ����V3�;�|";d�s�ȃ�k�8��������@u$�����0�і��VVVVV� 	   �p�������^Ë ^�jh���&����}��������k�84����E�   3�9^u6j
�����Y�]�9^uh�  �FP�F  YY��u�]��F�E������0   9]�t������k�8�����D8P�� �E������3ۋ}j
����YËD$�ȃ�k�8�������DP�� �jh��d����M��3��}�j����Y��u����g  j�<���Y�}��}؃�@�A  �4�������   �u�����   ;���   �Fu\�~ u9j
�����Y3�C�]��~ uh�  �FP�E  YY��u�]���F�e� �(   �}� u�^S�� �FtS�� ��8낋}؋u�j
����YÃ}� u��F����+����j8Y��������E�}��uyG�&���j8j �Bh��YY�E���ta������d� ���   ;�s�@ ���@
�` ��8�E������}�����σ�k�8�����DW�����Y��u�M���E������	   �E�� ����j�����Y�U����  ��f9E��   S�u�M��1���M�Q3�;�u�E�H�f��w�� ���]�   f9Es)�E�Pj�u�$  �����Et9�M싉�   f����q�M�jQj�MQPR�E�P�  �� ���Et�E�8]�t�M�ap�[��V�t$W3�;�u薓��WWWWW�    �5������   �F����   �@��   �t�� �F��   ��f��Fu	V�W  Y��F��v�vV�1��YP�i  ��;ǉF��   ���t�F�uOV��0�����Yt.V��0�����Yt"V��0����V�<�����0����k�8YY���)�@$�<�u�N    �~   u�F�tf� u�F   ��N�A���������	F�~���_^�U����UV�uj�X;��E�U�u�{����  �`���� 	   ����  S3�;�|;5d�r'�Q�����7���SSSSS� 	   ����������R  �ƃ�k�8��W�<����ƊH��u���������� 	   �j�����wP;Ӊ]��	  ���   9]t7�@$����E���HjYtHu���Шt����U�E�E��   ���Шu!蟑���腑���    SSSSS�$�����4����;��Mr�E�u�d��;�Y�E�u�M����    �U����    ����i  jSS�u�  ��D(�E���T,���AHtt�I��
tl9]tg��@�M8]��E�   �D
tN��L%��
tC9]t>��@�M�}��E�   �D%
u$��L&��
t9]t��@�M�E�   �D&
S�M�Q�uP��4�X ���|  �M�;��q  ;M�h  �M��D� ���  �}��  ;�t�M�9
u��� ��]�E��;؉]�E���   �M�<��   <t�CA�M�   �E�H;�s�A�8
u
AA�M�
�u�E�m�Ej �E�Pj�E�P��4�X ��u
�D ��uE�}� t?��DHt�}�
t����M��L�%;]�u�}�
t�jj�j��u��  ���}�
t�C�E�9E�G������D� @u����C��+E�}��E���   ����   K���xC�   3�@�����;]�rK�@���- t������-��u������ *   �zA;�u��@���AHt$C���Q|	���T%C��u	���T&C+���ؙjRP�u�  ���E�+]���P�uS�u�j h��  �� ���E�u4�D P蝎��Y�M���E�;EtP���Y�E�����  �E��  �E��3�;�����E��L0��;�t�M�f�9
u��� ��]�E��;؉]�E��   �E�f����   f��tf�CC@@�E�   �M����;�s!�Hf�9
u���Ef�
 �   �M�   �Ej �E�Pj�E�P��4�X ��u
�D ��uZ�}� tT��DHt'f�}�
t�f� ��M��L��M��L%��D&
�);]�uf�}�
t�jj�j��u�  ��f�}�
tf� CC�E�9E�������t�@u��f� f�CC+]�]������D j^;�u������ 	   ������0�h�����m�X����]��[���3�_[^��jh8��7����E���u������  襌��� 	   ����   3�;�|;d�r!藌���8�}���� 	   WWWWW������ɋ�����������k�8��L1��t�����;M�Au�I����8�/����    �P�l���Y�}���D0t�u�u�u�������E�������� 	   �����8�M���E������	   �E�薴����u����Yø�.á@���Vj^u�   �;�}�ƣ@�jP�_����YY�,�ujV�5@���^����YY�,�ujX^�3ҹ�.��,���� ����X1|�j�^3ҹ�.W����k�8������������t;�t��u�1�� B��H/|�_3�^��j<���=�� t�E���5,��&��Y�V�t$��.;�r"��81w��+�����Q�E����N �  Y^Ã� V�� ^ËD$��}��P�����D$�H �  YËD$�� P�� ËD$��.;�r=81w�`���+�����P� ���YÃ� P�� ËL$���D$}�`�����Q�ֵ��YÃ� P�� �U���SV�u�M��t'���u�3�9^u�u�u�]  YY�   �M;�u(����SSSSS�    �����8]�t�E��`p�3��h9]t�8tKW�E�(����D7t:u�P:Qt�P8t���:t@8u�8u��D0tA8tA8u�_����#�8]�t�M��ap�^[��j �t$�t$�'�����������7   ���"�.   ��������2��ƅp��������������
�t����
�t�����������������������ݽ`������a���u2����X銆�����-�&���
�t����
�t�������
�t�������`����؊�� ������k�����������U�������$�~$�   ��fD$f�f(�hf(5phf(�hf(�hf��%�  ��@  +�-�<  Ё�   ��(  fY�fX�f(�f\�fY�f(%�hfY�f(-�hf\�f~��ȃ�?������f\�f(��hfY�f(�fY�fX��Y��X�f�fo5Phf��fo5`hf��fs�.fY��X�fV�f��X���~  ��|  w�Y��X�fD$�D$��Ã���|$f�T$f�� f�$�,$����+�fo5@hf���  fn�fs�4fV���  fn�fs�4f$�$ft$�D$����f$$�$���$f$�l$��f�����  ���  s'�� t)�Z��   �r��+#��rJw�T$���9��r<��   ��   ��fD$�T$�ԃ��T$���T$�$����fD$����fD$�D$���=  �s1�D$=   �sfm�Y��   �fm�Y��   뉋T$=  �w�� u�D$=  �u� m��mú�  �V����D$%���=  �@s�fD$�X�l��fD$�D$��ÍI U�������$�~$�   ��fD$f��f%�f- 8f=���  f�f(0�fY��-�f(@�fX�f(P�f\�f-���� ) f(%`�fYك��Y��fY���f\�fYp������X�f(�f\�f5�����0mfT-��f(��f\�f��^�f\�f(x�\�fY�f\�f(H0fY�f(``fY��X�f(�fY�fX8fXH fY�fX`PfX�f(HpfY�fY�fX�f(H@fY�fX�f(�fY��Y�fY��   fY���fX����Y�f��X�f��X��\��X���f��   f��X��   �Y��X��   �X��X�f=���Y�f��   fT��Y��Y��   �\��\��   �\��Y����\��X��\��X��\ǃ��X�fD$�D$���?��f��f=~u���Y��f���Y��X��Y��f\$�D$����+������$        U����  3ŉE�SV�5<!3�9�W��u6SSjh$hh   S�օ�t��   ��D ��xu
��   9]~�M�EIf9t	@@;�u������+�E����u�u�u�u�u�u�u���  ��t;�uR9]�]�u��@�E9] u��@�E �u�rV  9E Yt���t�E �5� SSSS�u�uS�u �֋�;��}�u3��M  ~Bj�3�X����r6�G=   w�A)����;�t� ��  �P���;�Yt	� ��  ���E���]�9]�t�SSW�u��u�uS�u �օ���   SSW�u��=8!�u�u�׋�;���   ~?j�3�X����r3�F=   w�(����;�t� ��  �P�/��;�Yt	� ��  ���؅�txVS�u��u��u�u�ׅ�t]f�E t4�E3�;ǉu�tI;��p�VSP�u�tC  ����t0WWWWW�������!3�9EuPP��u�uVSj�u �� �E�S��6��Y�u���6���E�Y�e�_^[�M�3�������U����u�M��d���u$�M��u �u�u�u�u�u�q������}� t�M��ap���U���f�}��u�e� �bf�} s�E��3f�Af#E���E��@�u�M������E��p�p�E�Pj�EP�E�jP�]X  ����u!E��}� t�E�`p��E��M#���jhX��Ũ��3�3��}�j賬��Y�]�3��u�;5@���   �,���9tV� �@��uFf��xA�F���w�FP谫��Y����   �,��4�V�-���YY�,����@�tPV�z���YYF듋��b��j8��R��Y�,���,��9tFh�  � �� P��/  YY���,�u�4���Y�,������ P�� �,��<�}�;�t�g �  �_�_��_�O��E������   ������Ë}�j�Ǫ��Y��SVW�T$�D$�L$URPQQhԒd�5    �  3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�27  �   �C�D7  �d�    ��_^[ËL$�A   �   t3�D$�H3�����U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�6  3�3�3�3�3���U��SVWj j h{�Q�w�  _^[]�U�l$RQ�t$������]� U����$�S3�V�u�E��]�]��]��F�> t��<at9<rt,<wt�}��SSSSS�    �6�����3��I  �E  ��M��]��E	  �M�3�AF�:�W��  �Q� @  ;��+  ����S��   ��   �� �  ��tVHtG��t/��
t"���z  9]���   �M�E�   ��   	U��   �E@��   �M@�   �E�   �   �E��   �E������E�E����E��   9]�ut�M �E�   �r��TtZ��tDHt0��t����   f�E �uD	}�J9]�u:�e������E�   �59]�u%	}��E�   �$f�E �u�M �  �f�E t3���M   F�:������9]�tw�F�> t�jVh���]  ����ud��h�V��.  ��YYu���M   �;h�V��.  ��YYu���M   �h(�V�.  ��YYu���M   �F�> t�8t�{��SSSSS�    �+������h�  �u�E��u�uP�[  ����t3�� �E���M��H�M��X��X�X�H_^[��V�t$WV��������YtM�����u�@tu��u�@<tj�����j�������;�YYtV�����YP�� ��u
�D ���3�V�"����ƃ�k�8��������Y�D0 tW��z��Y����3�_^�jhx������E���u�z���  �{z��� 	   ����   3�;�|;d�r!�mz���8�Sz��� 	   WWWWW��������ɋ�����������k�8��L1��t�P�c���Y�}���D0t�u�����Y�E����y��� 	   �M���E������	   �E�蜢����u����Y�V�t$�F��t�t�v��	���f����3�Y��F�F^�U��QQ�EV�u�E��EWV�E��a������;�Yu�zy��� 	   �ǋ��J�u�M�Q�u�P�� ;ǉE�u�D ��t	P�ly��Y�ϋƃ�k�8�������D0� ��E��U�_^��jh��葡������u܉u��E���u�y���  ��x��� 	   �Ƌ���   3�;�|;d�r!��x���8��x��� 	   WWWWW�l������ȋ�����������k�8��L1��u&�x���8�x��� 	   WWWWW�+�����������[P����Y�}���D0t�u�u�u�u�������E܉U���>x��� 	   �Fx���8�M���M���E������   �E܋U��Ԡ����u�����Y�U��$������  �  3ŉ�  ��$  V3�9�(  �E��u��u�u3��t  ;�u'��w���0�w��VVVVV�    �Z���������I  ��   S�ރ�k�8����W�<����ÊH$������}��M�t��u3��(  ����u&�jw��3��0�Nw��VVVVV�    ���������  �@ tjj j V������V�%;  ��Y��  ��D���  �:b���@l3�9H�E���P��4��� !����  ��t
�}� ��  �� �e� ��(   �u��E��u���  �e� ��u��E����  �3�<
����P�M�������Yuj�E�VP�0Z  �������  �0�E�+��(  ����  j�E�VP�Z  �������  F�E�3�PPj��  Qj�M�QP�u�F�E��u��� �����O  j �E�PV��  P��4�� ���%  �E�E�;��   �}� ��   j �E�Pj��  P�ƅ  �4�� ����  �}���  �E��E��d<t<u�3�f��
��FF�E��M��u��U�<t<u9�u��HW  f;E�Y��  �E��}� tjXP�E��(W  f;E�Y�t  �E��E���(  9E��y����c  ���@��%  �E�3��}� �u���   9�(  �E��e  �M��e� +M��E�;�(  s'�U��E��A��
u
�E�� @�E��@�E��}�   rы��E�+�j �E�PV�E�P��4�� ����  �E�E�;���  �E�+E�;�(  r��  �}���   9�(  �E���  �M�3�+M��E�;�(  s1�U��E��AAf��
u�E�f�  @@FF�}�f�@@FF���  rǋ��E�+�j �E�PV�E�P��4�� ���'  �E�E�;��"  �E�+E�;�(  �w����  9�(  �E��-  �M��e� +M�j���  ^;�(  s,�U��u��f��
u
f�  �u�u�f�Ɓ}�R  r�3�VVh�  ��  Q���  +��+���P��PVh��  �� ��;�tyj �E�P��+�P��5  P�E�� �4�� ��t	u�;���	�D �E�;�G�E�+E�;�(  �E��6����0j �M�Q��(  �u��0�� ��t�E��e� �E��	�D �E��E���uV�}�3�9u�t j^9u�u�r��� 	   �+�u��r��Y�'��D@t�E��8u3���nr���    �vr���0����+E�_[��  3�^�������  ��jh��貚���E���u�;r���  � r��� 	   ����   3�;�|;d�r!�r���8��q��� 	   WWWWW�������ɋ�����������k�8��L1��t�P����Y�}���D0t�u�u�u�������E���q��� 	   �q���8�M���E������	   �E��2�����u�R���Y�jh���֙���E���u�Lq��� 	   ����   3�;�|;d�r�+q��� 	   SSSSS��������Ћ����<�������k�8��L��t�P�;���Y�]���Dt1�u����YP�!��u�D �E���]�9]�t��p���M��p��� 	   �M���E������	   �E��Q�����u�q���Y��������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��V�t$V��������Yu� p��� 	   ���^�W�t$j �t$P�� �����u�D �3���tP��o��Y�����ƃ�k�8�������D0� ���_^�jh�������E���u�o���  �o��� 	   ����   3�;�|;d�r!�uo���8�[o��� 	   WWWWW��������ɋ�����������k�8��L1��t�P�k���Y�}���D0t�u�u�u��������E����n��� 	   � o���8�M���E������	   �E�蕗����u����Y�U���SW�}3�;�u �n��SSSSS�    �Q���������c  W�r��9_Y�E�}�_jSP�������;ÉE�|ӋWf��u+G�,  ��OV��+����u�tA�u��U���k�8�������D2�t��;�s���:
u�E�3�B;�r�9]�u�E���   ��x��n���    �   �G��   �W;�u�]��   �u��]���k�8+���������E��D0�twjj �u��
�����;E�u�G�M��	�8
u�E@;�r�f�G  �?j �u��u����������}����9�   9Ew�O��tf�� t�G�E��D0t�E�E)E��E�M��^_[���@@t�x tP�t$��P  f=��YYu�����U��V����u�E�M������>�Yt�} �^]��G@SV����t9� u3�D$�2��L$P������CC�>�Yu�l���8*uj?���r���Y�|$ �^[�U��$�����t  �  3ŉ��  ���  S��  V��   W��  3��M��Eĉ]؉}��}�}ȉ}�}Љ}��}��	��9}�u-�2l��WWWW�    W��������}� t�E��`p�����K  ;�t��3�f;׉}ԉ}��}��U��  j_��}� �u��  �B�f=X w��������3�����j��Y;��E���  �$���3��M���E��E��EȉEЉE�E��  �� t>��t-��t+�t���c  �M��Z  �M��Q  �M��H  �M�   �<  	}��4  f��*u ���]؋[��ۉ]��  �M��]��  �E�k�
�ʍDЉE���  �e� ��  f��*u���]؋[��ۉ]���  �M����  �E�k�
�ʍDЉE��  ��ItH��ht:��lt��w��  �M�   �  f�>lu��M�   �u��z  �M��q  �M� �h  �f=6 uf�~4u���M� �  �u��F  f=3 uf�~2u���e�����u��'  f=d �  f=i �  f=o �	  f=u ��  f=x ��  f=X ��  �e� �E�R�u��E�   ������  ��d��  �   ��S��   t_��At+�tA+�t+���  �� �E�   �U܃M�@�}� �u�   �u�E���  �E�   �<  f�E�0��   �M� �   f�E�0u�M� �}���u�������E� �]؋[��]���  ��u�|)�E�e� ���u���  �����  �M���QP�������YYtFF�E�9}�|���  ��X�C  +�tg+��8���+���  ���3�F�E� �ủ]؉E�t-�E��E�P�E��E� ���   �E�P�E�P�1K  ����}	�u��f�E��E��E�u��M  ������]�t-�H��t&f�E� � �M�t�+��E�   �  �e� �  �|)�E�P�|3��Y��  ��p��  �u  ��e��  ��g�k�����itY��nt��o��  �E��E�   tI�M�   �@�3���]��#������  �E� t	f�E�f���Eԉ�E�   �  �M�@�E�
   f�E� ��D  ��S���p  uf��guE�E�   �<9E�~�E�}�   ~+�}��]  W�o:�����U�Y�E�t
�E�}�����E�   ����E��C��E��E�P�u����u�]�P�u��E�VP�5�&�P��Y�Ћ]����   t�}� u�E�PV�5�&��O��Y��YYf�}�gu��u�E�PV�5�&��O��Y��YY�>-u�M�   F�u�V�q����E�   �M��!��s�<���+���������V  �E�'   �E��E�   ������E���Qf�E�0 f�E��}�����f�E� ��������E� t�E�@�]�t�C���C����E�@�C�t��3҉]��E�@t��|��s�؃� �ځM�   f�E� ��ڋ�u3ۃ}� }	�E�   ��e���   9E�~�E���u!EЍ��  �E��M�����t$�EܙRPSW�x+  ��0��9�]�����~M��N�̍��  +�Ff�E� �E��u�tD��t�΀90t9�M�M��0@�*��u��)�E�E��E�   �	Of�8 t@@��u�+E����E��}� ��   �E�@t+f� tf�E�- ��tf�E�+ �
�tf�E�  �E�   �]ȋu�+�+]��E�u�učE�Sj �������uЋ}čEԍM�������E�Yt�E�uWSj0�E��������}� uN��~J�}�u��M܍E�P�E����   �E�WP�G  �����E�~�u��Eču�� ���}��}� Y���M����M�V�E��L���Y�}� |�E�t�učE�Sj �������}� t�u��8����e� Y�u��f���E�t$�M��]؋��������c���    3�PPPPP�����}� t�E��`p��Eԋ��  _^3�[�B������  ���ǥ�2�m�v�����V�t$V�]��P�'  ��YYt{������ ;�u3��������@;�u_3�@��f�FuNSW�<���? �   u S�P6����Y�u�Fj�F�X�F�F��?�~�>�^�^�N  _3�[@^�3�^Ã|$ t'V�t$f�F tV����f�����f �& �f Y^������������WVS3��D$�}G�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u�L$�D$3���؋D$����A�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�Ou���؃� [^_� QV��L������u��a���    3��)�~D u j$�
5����Y�FDu��a���    �D$��FD^Y�U��SVWj j ��	  ���  V�5 2����	  �}����f%�f=�QQ��   �02�}��E�$�  ��YY~O��~"��uE�ESQ��EQ�$j�i  ���   �E����E�\$���$�;$  �]VS�b	  ���]�ES��$����\$�E�$jj�j  ���9�E�$��#  �E�Y�mY�]���]����Dz	f�� �f	}VS�	  YY�E_^[]�U��QQSV���  V�5$2��  �EYY�؋EQf%�f=�Q�$uU��   ��YY~-��~��u#�ESQQ�$j�~  ���rVS�  �EYY�d�ES��$���\$�E�$jj�?�+#  �]��EY�]�Y����DzVS�T  �E�YY�"�� u��E�S���\$�E�$jj�]  ��^[��U��QQ�E�E�M�]��  ��������f�E��E���U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]ËM��  #�f;�uj��f���u�E�� u9Utj��3�]�U�����U����Dz3��   3�f�E�uc�E�� u9MtU�]��������Au3�@�3���e�E   �t�M�eJ�Et�f�e��;�tf�M ��EQQQ�$��������%Q���EQQ�$������U�����  �����  �E�]�U��E�MSVW3��x�E3ۉx�EC���xt�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H��  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP��  �EPSj �u�( �M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]�U��j �u�u�u�u�u�u�
�����]�U����ESV3ۋ���C��u�t�]tS��  Y����  �t�Etj��  Y����w  ����   �E��   j�  �EY�   #�tT=   t7=   t;�ub��M����82��{L�H��M�����{,�82�2��M�����z�82���M�����z�(2��(2��������   ���   �E��   3��t����W�}�����D��   ��E�PQQ�$�/����M��]��� �����������}�E�����$�T���]�����Au���3��E�����f�E�����;�}"+��]�t��u���m��]�t�M�   ��m�Hu���t�E����]��E������_tj�h  Y�e���u��Et�E tj �M  Y���3���^��[�ËD$��t~����Y��� "   ��Y��� !   ÊD$� tj��t3�@ètj��tjX�������U��� 3���P2;Mtd@��|�3����E�t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E��g  �E�P��)  ����uV�:���Y�E�^�Ë�T2�h��  �u(�4  �u�����E ����U��=�3 u(�u�E���\$���\$�E�$�uj�3�����$]��X��h��  �u� !   ��   �EYY]�U������   �  3ĉD$|�u �EP�u��������u%�d$@�P�EP�EP�u�E �uP�D$P�������u�������=�3 u+��t'�u �E���\$���\$�E�$�uP������$�P�#����$��  �u �+   �EYY�L$|3��q�����]�Q��<$�$Y�Q�<$���$Y�U��Q��}��E�M#M��#E�����E�m�E���QQ�L$��t�-83�\$���t����-83�$������t
�-D3�$���t	�������؛�� t���$�YY�jh����3�9��tV�E@tH9P3t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%P3 �e��U�E�������e��U�����������������ƅp�����   
�t{��   ���N�����-`3�ٛݽ`������a���Aud�m   
�t[���   ���   �����ƅp�����J   
�t3�r   ���������TS�����- )�T�����- )���h����S���wh��ƅp����7S��������3��{h������a���t	�(   ������@u����������R���   ��
�u�����������
�u�������������U�������$�~$�   ��fD$�    f(�f�fs�4f�� f(��f(��f( �f(%Єf(5��fT�fV�fX�f�� %�  f(���f(���fT�f\�fY�f\��X�fY�f(�fXƁ��  �����  ��   ���  ��*�f���
��   �    �� D�f(p�f(�f(��fY�fY�fX�f(���Y�f(-��fY�f(� �fT�fX�fX�fY��Y�fX�f(��fY�f(�f�fY˃�f(�fX�f��X��X��X�fD$�D$���fD$f(0���� f�� �� wH���t^���  wlfD$f(��f( �fT�fV���� f�� �� t�X�ú�  �Of ��^�fP��   �4f@��Y���������������  ���  s:fW��^ɺ	   ��fL$�T$�ԃ��T$���T$�$詙���D$���fT$fD$f~�fs� f~с��� ��� t���  릍�$        �L$f�9MZt3�ËA<��8PE  u�3�f�x�����������̋D$�H<��ASV�q3҅�W�Dv�|$�H;�r	�X�;�r����(;�r�3�_^[���������������U��j�h8�h@:d�    P��SVW�  1E�3�P�E�d�    �e��E�    h   �<�������tU�E-   Ph   �R�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]ËD$�����������ËD$�L*V9Pt��k�t$��;�r�k�L$^;�s9Pt3���5����:��Y�j hX��z��3��}�}؋]��Lt��jY+�t"+�t+�td+�uD�-<�����}؅�u����a  �����`�w\���`���������Z�Ã�t<��t+Ht�&Q���    3�PPPPP�������뮾�������������
�������E�   P��9���E�Y3��}���   9E�uj���9E�tP�2}��Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.�@*�M܋D*�@*�9M�}�M�k��W\�D�E����f9����E������   ��u�wdS�U�Y��]�}؃}� tj ��{��Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3��x��ËD$��ËD$����t$�!3�@� jhx��?x��3��}��5���8��Y��;�uS�E�P���Y;�tWWWWW�F������}�t!h���h ;�thЍP�d ��;�u���V�8��Y���}��u�u�։E��/�E� � �E�3�=  �����Ëe�}�  �uj�� �e� �E������E���w���U���V�u�M��V����U3�;�u/��N��VVVVV�    �������}� t�E�`p�������  S�];�u/�N��VVVVV�    �Q������}� t�E�`p������  �E�9pu$�E�PSR������}� �u  �M�ap��i  W�   f�
����B�D�UtY�: u3��lj�p�M�jQjJRW�p�E�P軴����$��uf�E������   f�E�f�M�f��f��E���E���э�Atf��  �����f�����C�DtU�; u3��hj�p�M�jQj�K�QW�p�E�P�2�����$��uf�E����uHf�E�f�M�f��f��ȋE�C��э�Atf��  �����f;�u,f��t<�U������2M���    �}� t�E�`p������$���H�}� t�M�ap���}� t�E�`p�3�_[^��j �t$�t$��������j �t$�t$�t$�t$�v2  ���S�\$U3�;�u3��=VWS�����FV������;�YYt SVW��<������tUUUUU�2��������3�_^][�U���S�u�M�����3�9]u.�SL��SSSSS�    �������8]�t�E�`p������   V�u;�u.�L��SSSSS�    ������8]�t�E�`p������   W�}�9_uV�u�'��YY�{�Ef�����@�D:�Et� :�u3��3��E�����f�����F�D:t�:ӈU�u3��3Ҋ�F�U���f;�uf;�u�8]�t�E�`p�3�_^[�����H8]�t��M�ap���j �t$�t$��������U���S3�9]u�/K��SSSSS�    �������3��jV�u;�u�K��SSSSS�    �������9ur3��>�u�M��A����M�9Y�F�tH9Ew
��D
u���+ȃ�+�N��8]�t�M��ap�^[��j �t$�t$�Z������U��QQ�  3ŉE���SV3�;�W��u:�E�P3�FVh$hV�!��t�5��4�D ��xu
jX���������   ;���   ����   9]�]�u��@�E�5� 3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w������;�t� ��  �P�)���;�Yt	� ��  ���؅�ti�?Pj S�������WS�u�uj�u�օ�t�uPS�u�!�E�S�&����E�Y�u3�9]u��@�E9]u��@�E�u�  ���Yu3��G;EtSS�MQ�uP�u�2  ����;�t܉u�u�u�u�u�u�!;��tV�'���Y�Ǎe�_^[�M�3��u�����U����u�M��.����u$�M��u �u�u�u�u�u�������}� t�M��ap���3�@�|$ u3��U��SVWUj j h���u�W  ]_^[��]ËL$�A   �   t2�D$�H�3������U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h��d�5    �  3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y��u�Q�R9Qu�   �SQ��3�SQ��3�L$�K�C�kUQPXY]Y[� ��������U��W�}3�������ك��E���8t3�����_��U����u�M��x����E����   ~�E�Pj�u�%���������   �M�H���}� t�M��ap��Ã=�� u�D$��-�A���j �t$����YY�U���(�  3ŉE�SV�uW�u�}�M�������E�P3�SSSSW�E�P�E�P��8  �E�E�VP�8.  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[������U���(�  3ŉE�SV�uW�u�}�M��G����E�P3�SSSSW�E�P�E�P�#8  �E�E�VP��2  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�������U��MSV�u3�;�W�yu�LE��j^�0SSSSS����������   9]v݋U;ӈ~���3�@9Ew�E��j"Y�����;��0�F~�:�t��G�j0Y�@J;��M;ӈ|�?5|�� 0H�89t�� �>1u�A��~W���@PWV�l�����3�_^[]�U��Q�U�BS��VW��% �  ��  #ωE�B��پ   �%�� �ۉu�t;�t�� <  �(��  �$3�;�u;�u�Ef�M�X��L��<  �]����������M��E���ΉH�u��P������Ɂ���  �։P�t�M�_^f�H[��U���0�  3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���u�����f��<  �uЉC�E։�EԉC�E�P�uV��3����$��t3�PPPPP�*������M�_�s^��3�[����������������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j���Y�U��E�M%����#�������Vt1W�}3�;�tVV�,E  YY��B��j_VVVVV�8��������_��u��P�ut	��D  ����D  YY3�^]�U������   �  3ĉ�$�   �E�SV�u�HW�L$t+Ht$HtHtHtHHtHutj��   �hj�
j�j�j[Q�~WS���������uG�E��t��t��t�d$P���L$P�F����\$@���L$PW�NQPS�D$P�D$$P�V�����h��  �t$�^����>YYt�=�3 uV��  ��Yu�6�%���Y��$�   _^[3�耻����]�jh���Zi���e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E��\i���U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�^�����t3�@�3�[���������3��U��� SVW�3)��3�9P��E��]��]�]���   hl��!��;��y  �5d h`�W��;��c  P�z(���$P�W�P���P�e(���$<�W�T���P�P(���X��E�P�����YYtSSSSS�>������}�u,h �W��P�(��;�Y�`�th�W��P�(��Y�\��\��M�;�ty9`�tqP�Z(���5`����M(��;�YY��tV;�tR��;�t�M�Qj�M�QjP�ׅ�t�E�u3�E�P�(����YtSSSSS蟼�����}�r	�M    �D�M   �;�T�;E�t1P��'��;�Yt&��;ÉE�t�X�;E�tP��'��;�Yt�u��ЉE��5P��'��;�Yt�u�u�u�u����3�_^[�ËD$S3�;�VWt�|$;�w�U>��j^�0SSSSS����������=�t$;�u��ً�8tBOu�;�t��
BF:�tOu�;�u��>��j"Y����3�_^[�U��SV�u3�9]Wu;�u9]u3�_^[]�;�t�};�w��=��j^�0SSSSS�n���������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x�����T=��j"Y���낋L$V3�;�|��~��u�h�^áh��h�^��=��VVVVV�    輻�������^�QQ�D$���$�$YY�U��QQ��E�]��E��E3E%���3E�E��E���U��E��  ��#�f;�u-�EQQ�$�����HYYtHtHt3�@]�j�jX]ø   ]�% �  f�ҋ�u�E�� u�} t�������   ]����]����D��z��������@]����%���   ]���h   �P����Y�L$�At�I�A   ��I�A�A�A   �A�a �ËD$���u��;��� 	   3��V3�;�|;d�r��;��VVVVV� 	   �j�����3�^Ëȃ�k�8�������D��@^�U���SV�u3�;�W�}u;�v�E;�t�3���E;�t�������v�[;��j^SSSSS�0����������R�u�M������E�9X��   f�Ef=� v6;�t;�vWSV�M������;��� *   �;��8]�� t�M��ap�_^[��;�t.;�w(��:��j"^SSSSS�0聹����8]�t��E��`p��u�����E;�t�    8]��0����E��`p��$����MQSWVj�MQS�]�p�� ;�t9]�b����M;�t����D ��z�H���;��k���;��c���WSV�z������S���j �t$�t$�t$�t$��������������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� �A@t�y t$�Ix��������QP�N��YY���u	���U��V����M�E�M�����>�t�} �^]��G@SV����t4� u.�D$�-��L$������C�>�u��8���8*u�ϰ?�i����|$ �^[�U��$�����x  �  3ŉ��  ��   S��  V3�W��  ��  �M��EЉ}ԉu��u�u��u��uĉu��u������9u�u-�|8��VVVV�    V�������}� t�E��`p������  �E��@@��   P�"������Yt6�u��������Yt(�u������u����4����������k�8YY3����)�@$�u����u���������Yt6�u���������Yt(�u������u����4���������k�8YY3����)�@$��"���;�������҉ủu؉u��u��U��  C3�9Ẻ]���  �ʀ� ��Xw����X����M�k�	��x�j��^;ƉE���  jY;��z  �$��3��M���E��E��E��EĉE�E��V  �� t<��t++�tHHt���8  	u��0  �M��'  �M��  �M�   �  �M��	  ��*u ���}ԋ����}���  �M��]���  �E�k�
�ʍDЉE���  �e� ��  ��*u���}ԋ����}���  �M���  �E�k�
�ʍDЉE��  ��ItF��ht8��lt��w�w  �M�   �k  �;luC�M�   �]��V  �M��M  �M� �D  �<6u�{4uCC�M� �  �]��'  <3u�{2uCC�e�����]��  <d�  <i��  <o��  <u��  <x��  <X��  �e� �e� �E�P��P�a���Y���E�Yt�MЍu�������C���]���  �MЍu�������  ��d�t  ��  ��S��   t[��AtHHtAHHtHH�K  �� �E�   �U�M�@�}� �]�   �]܉E���  �E�   �  f�E�0uu�M�   �lf�E�0u�M�   �M����u������f�E��}ԋ��}���  ��u��)�E܋E��E�   �  ��X�4  HHt]+��c���HH��  ��f�E��}�t'�G�Ph   �E�P�E�P��������t�E�   ��G��E��E�   �E�E��L  ������}�t/�H��t(f�E� � �M�t�+����E�   �  �e� �  �|)�E�P�,���Y��  ��p��  �r  ��e��  ��g�������itU��nt��o��  �E耉u�tI�M�   �@�7���}��m�������  �E� t	f�E�f���Ẻ�E�   �  �M�@�E�
   �M�f���A  ��G��W��i  u��guH�E�   �?9E�~�E��}�   ~.�u���]  V�$�����U�Y�E�jt
�E܉u�����E�   ^��G��E��G��E��E�P�u����u��}�P�u��E�SP�5�&����Y�Ћ}����   t�}� u�E�PS�5�&���Y��YY�}�gu��u�E�PS�5�&���Y��YY�;-u�M�   C�]�S�t����u��M��!��s�u���HH��������Z  �E�'   �E��E�   ������E�Q�E�0�E��E�   ����f�� ��������� t��@�}�t�G���G�����@�G�t��3҉}���@t��|��s�؃� �ځM�   f�E� ��ڋ�u3ۃ}� }	�E�   ��e���   9E�~�E����u!Eč��  �E��M������t$�EؙRPSW�4�����0��9�]�����~M��N�̍��  +�Ff�E� �E؉u�tM��t�΀90tB�M܋M��0@�3If�8 t@@��u�+E������u�|)�E܋E��I�8 t@��u�+E܉E؃}� ��   �E�@t%f� t�E�-��t�E�+��t�E� �E�   �]�+]�+]��E�u�uЍE�Sj �.������uċ}ЍE̍M��>����E�Yt�E�uWSj0�E��������}� �E�tQ��~M�u܉E���M�Pj���  P�E�FPF���������u9E�t�u��E̍��  ������}� Yu���M����M�P�E�����Y�}� |�E�tWSj �E��������}� t�u������e� Y�]�����E�t!�}Ԋ�� ����/���    3�PPPPP����3�9u�t
�}�������}� t�E��`p��E̋��  _^3�[�������  �Ð��<�Y������� ��3��V�t$����  �v�K����v�C����v�;����v�3����v�+����v�#����6�����v �����v$�����v(�����v,������v0������v4�����v�����v8�ܾ���v<�Ծ����@�v@�ɾ���vD������vH蹾���vL豾���vP詾���vT衾���vX虾���v\葾���v`艾���vd聾���vh�y����vl�q����vp�i����vt�a����vx�Y����v|�Q�����@���   �C������   �8������   �-������   �"������   �������   �������   �������   ��������   �������   �������   �ս����,^�V�t$��t5�;�4tP跽��Y�F;�4tP襽��Y�v;5�4tV蓽��Y^�V�t$��t~�F;�4tP�v���Y�F;�4tP�d���Y�F;�4tP�R���Y�F;�4tP�@���Y�F;�4tP�.���Y�F ;�4tP����Y�v$;5�4tV�
���Y^���������������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^��U����  3ŉE�j�E�Ph  �u�E� �!��u����
�E�P�  Y�M�3�腦����U���4�  3ŉE��E�M�E؋ES�EЋ V�E܋EW3�;E�M̉}��}��_  �5x �M�QP�օ��� t^�}�uX�E�P�u�օ�tK�}�uE�u܃���E�   u�u��������YF;�~[�����wS�D6=   w/�4�����;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P芺��;�Yt	� ��  ���E���}�9}�t؍6PW�u��,�����V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u�� ��t`�]��[9}ԋ� uWWWWV�u�W�u�Ӌ�;�t<Vj�����;�YY�E�t+WWVPV�u�W�u��;�u�u�蟺��Y�}���}��t�MЉ�u�����Y�E��e�_^[�M�3��Ӥ����U����  3ŉE��}�SVW}3���  � ��5!3�3�C;�u3�E�PSh$hS�օ�t� ���D ��xu
jX� ��� �;�u�u�u�u�u���  ��t;�u�9} �}�u�E� �@�E 9}u�E� �@�E�u �U���9EYt���t�E�� WWWW�u�uW�u�Ӌ�;��u��6���~;���w6�F=   w�.�����;�t� ��  �P蠸��;�Yt	� ��  ���E���}�9}������VW�u��A�����WWV�u��u�uW�u�Ӆ���   �F;�~D=���w=�D6
=   w������;���   ���  ���P�!���;�Yt	� ��  �����3�;�tb9} u�E� �@�E �}S�u���u��4�uf����u f�N����!f�~����E�tf�>��uWS�u��������e� S�����Y�u�������E�Y�e�_^[�M�3�询����U����u�M��h����u �E��u�u�u�u�uP�������}� t�M��ap���U���4S3��E�VW���]܉]؈]��E�   �]�t	�]��E��
�E�   �]��E�P�h2  ��YtSSSSS�>������E�P�u�����YtSSSSS�#������M� �  ��u�� @ u9E�t�M������+ú   ��   �tGHt.Ht&�E'������('��j^SSSSS�0�ȥ������  �U����t��   u��E�   @��}��EjY+�t7+�t*+�t+�t��@u�9}����E���E�   ��E�   ��E�   ��]��E�   #¹   ;��   ;t0;�t,;�t=   ��   =   �@����E�   �/�E�   �&�E�   �=   t=   te;������E�   �E���E�   t�t���#M��x�E�   �@t�M�   �M�   �}�u�M�f� t	}�� t�M�   ��E�   롨t�M�   �ݏ������u��%������%���    �   �E�=!S�u��    �u�E�P�u��u��u�׃���E�um�M��   �#�;�u+�Et%�e����S�u�E��u�P�u��u��u�׃���E�u4�6�ƃ�k�8�������D0� ��D P�H%��Y�%��� �  �u��H ;�uD�6�ƃ�k�8�������D0� ��D ��V�%��Y�u��� ;�u���$���    룃�u�M�@�	��u�M��u��6肌����Ѓ�k�8������YY�M����L��Ѓ�k�8�������D$� ��M��e�H�M���   ����G  �Etqj���W�6�)�����;ǉE�u�C$���8�   tM�6���������j�E�P�6�]�腑������u�}�u�E�RP�6�P,  ��;�t�SS�6�̳����;�t��E����   � @ �M� @  u�E�#�u	}�	E�E#�;�tD=   t)= @ t"=   t)= @ t"=   t= @ u�E���M�  #�;�u	�E���]��E   tO�E�@�]�uF�E��   �#�=   @��  =   ��G  ;�u"�E�;�v���  ����   ���  ��ȃ�k�8�������D$�2M���0��ȃ�k�8�������D$�M�������
�8]��u!�Et��ȃ�k�8�������D� �}��   ���#�;���  �E��  �u��� S�u�E�jP�u������W�u�!�����  �D P�f"����ȃ�k�8�������D� ��6�w���Y�����jSS�6�j��������   SSS�6�U���#���������j�E�P�6�V���������������tg����   �}�﻿ uU�E������E�;����������   �������jSS�6�������tySSS�6�է����#���_����=����E�%��  =��  u�6����Y�I!��j^�0���   =��  uSj�6���������������E�����SS�6���������E�3�HtH������E���  �E�   ��E�﻿ �E�   �E�+�P�D=�P�6舮�������t�9}�������6�~���Y� ��� �E���6����������k�8���_^[��jh����H��3��u�3��};���;�u�_ ��j_�8VVVVV����������Y��3�9u��;�t�9ut�E%������@tu��u�u�u�u�E�P���0������E��E������   �E�;�t���H���3��}9u�t(9u�t�������k�8�����D� ��7褉��Y�U��j�u�u�u�u�u������]�U���S3�9]u3��=  W�u�M��׼���}�9_u&�u�u�u�'�����8]��  �M��ap��  9]u.�@��SSSSS�    �ߝ����8]�t�E��`p�������   V�u;�u.�
��SSSSS�    詝����8]�t�E��`p������   �Ef��M����@�D:�Et,9]u�3��D8u^���F� :�u3��3��E�����f�����F�D:t9]u3����M:�t�3ۊ�F����3�f;�u!f;�t	9]�v���8]�t�E��`p�3�^_[�����H8]�t��M��ap���j �t$�t$�t$�������U����  3ŉE�V3�95�5tN�=�5�u��(  ��5���uf���pV�M�Qj�MQP�(!��ug�=�5u��D ��xuЉ5�5VVj�E�Pj�EPV�$!P�� ��5���t�V�U�RP�E�PQ� !��t�f�E�M�3�^���������5   ��U���SV�u3�;�t9]t8u�E;�tf�3�^[���u�M�聺���E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P�Ѓ����YYt}�E����   ��~%9M| 3�9]��R�uQVj	�p�� ���E�u�M;��   r 8^t8]����   �e����M��ap��Y������� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p�� ���:����j �t$�t$�t$��������U����  3ŉE�SV�u�F@W��  V�������Y��)t.V�׹�����Yt"V�˹����V����軹����k�8YY��Ǌ@$$<�A  V蚹�����Yt.V莹�����Yt"V肹����V�����r�����k�8YY��Ǌ@$$<u\�N�]x����A����VP�0��YY���u	f����   �Nx��8��A����VP��/��YY���t�f����   V��������Yt.V�������Yt"V������V�����Ѹ����k�8YY����@�t^�u�E�jP�E�P���������l���3�9]�~4�Nx��L���A���D�VP�G/��YY����7���C;]�|�f�E� �F�x��Ef����EVP�%  YY�M�_^3�[������U���S3�9]V�uu;�u9]u3���  ;�t9]w���j^SSSSS�0还��������  9]u���W�};�u�����j^SSSSS�0莘�����(  �u�M��+����E�9Xu�uW�uV�������L  �}��U��u��@G:�tJu����@G:�tJt�Mu�9]u�@;���   8t�}u5�x�;��}�r�E�P�E�� P�������YYt�M�9u�s��+E����   �}�uZ�E��v:�|�;��}r!�E�P�E� P������YYt�M9us�E��+M��t���\�8]�t�E�`p�jPX�   �����j"^SSSSS�0�m�����8]�t�E�`p����d��+΃�|M�x�;��}r�E�P�E� P�"�����YYt�M9us��+E�t��j����j*X�8]�t�M�ap��8]�t�E�`p�3�_^[��j
j �t$�j   ���U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  �������W�M�E�u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5�5N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r;�ur��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC��5��+�5;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5�5N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3���5A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;�5��5��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}硤5��5�3�@�   ��5�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+�5��M���Ɂ�   �ً�5]���@u�M�U�Y��
�� u�M�_[��U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  �������W�M�E�u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5�5N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r;�ur��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC��5��+�5;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5�5N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3���5A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;�5��5��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}硼5��5�3�@�   ��5�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+�5��M���Ɂ�   �ً�5]���@u�M�U�Y��
�� u�M�_[��U���|�  3ŉE��ES3�V3��E��EF3�9]$W�E��}��]��u��]��]��]��]��]��]��]�u�_��SSSSS�    �������3��  �U�U��< t<	t<
t<uB��0�B���/  �$�J
�Ȁ�1��wjYJ�݋M$�	���   �	:ujY������+tHHt����  ���jY�E� �  뢃e� jY뙊Ȁ�1���u�v��M$�	���   �	:uj�<+t(<-t$:�t�<C�<  <E~<c�0  <e�(  j�Jj�y����Ȁ�1���R����M$�	���   �	:�T���:��f����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�]���<+t�<-t��`����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*�<	�u��n���j�����J��M��Ȁ�1��wj	��������+t HHt���;���j�����M��jY�@���j�o����u���B:�t�,1<v�J�(�Ȁ�1��v�:�뽃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�[����B:�}��O����M��E�O�? t�E�P�u��E�P�@  �E�3Ƀ�9M�}��E�9M�uE9M�u+E=P  ��  =������  ��5��`;��E���  }�ؾ@7�E���`9Muf�M�9M���  �E��}���T�����u��q  k�Ƌ�f�; ��]�r��}�����M��u��]��]��S
�M�3��E��EԉE؉E܋¿�  3�#�#�% �  f����<
����  f�����  f������  f���?w3��EȉE���  f��uG�E����u�}� u�}� u	f!M���  3�f;�u!G�C���u9Ku9u�M̉MȉM��  !M��u��E�   �M��U�Ʌ҉U�~U�Lă��M��]��M��U���	�e� �ʋV��
;�r;�s�E�   �}� �^�tf��E��m��M��}� ��]�FF�E��M��}� ����  f��~;�E�   �u-�u؋M��e�������M����ʁ���  f���u؉M��f��M����  f��}B��������E�t�E��M܋]؋U��m�����ًM������N�]؉M�u�9u�tf�M�f�}� �w�Mԁ��� �� � u3�}��u*�e� �}��u�e� f�}���u	f�E� �G�f�E���E���E�f����u�sf�M�f�MċM؉MƋM���M�f�}��f����e� %   � ���e� �Ẽ}� �m����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W�M�_^3�[貁����R��/t���z)U���t�  3ŉE�S�]VW�u�}�f��U��ʸ �  #ȁ��  f�ɉ]��E���E���E���E���E���E���E���E���E���E���E���E�?�E�   �M�t�C-��C f�ҋu�}�u.��u*��u&f!;f;�����$ �C�C�C0�C 3�@��  f�����   �   �;�f� u��t��   @uhĶ�Qf��t��   �u��u;h���;�u0��u,h���CjP�#�����3���tVVVVV�z������C�*h���CjP�������3���tVVVVV�N������C3��  �ʋ�i�M  �������Ck�M���������ىM�3���5�ۃ�`;�f�U�u�}�f�E��M���  }�@7�ۃ�`�M�;���  �E�T�˃������y  k�M�f�9 ��M�r��}ĥ��Eĥ�MƉE����y
�U�3��Ͼ�  3�#�#��E��E��E�E��� �  f;֍���  f;���  f=����  f=�?w3��E�E�E���  3�f;�u@�E����u9u�u9u�u	f�u���  f;�u$�U�@�B���u9ru92u�u�u�u��  �}�u��}��E�   �U��u�҅��u�~X�T��U��U����U��U��u��6����փe� �4;�r;�s�E�   �}� �}��w�tf��E��m��M��}� �GG�E��M��}� �}���  f��~;�E�   �u-�U��}�u��e������U�������  f���}�U��f��R��  f��}H�����҉U���E�t�E��U��}�u��m�������U�������M��}�U�uσ}� tf�M�f�}� �w�U����� �� � u3�}��u*�e� �}��u�e� f�}���u	f�E� �@�f�E���E���E�f=�sf�U�f�U��U�U�U���U�f�E��f��Ƀe� ��   ��� ���e� �M���k���3��M���f���?��  �H  �u��E��ы�3�#�#�� �  f;Ӎ<�E��E��E�E�����  f;���  f������  f���?w�E���  f;�uG�E����u9E�u9E�u	f�E���  f;�uG�E����u
9E�u9E�t��e� �E��E�   �U��u�҅��u�~R�u؍T��u��U��U��u��6��e� �֋p��;�r;�s�E�   �}� �X�tf� �E��m��M��}� �@@�E��M��}� ����  3�f;�~<�E�   �u.�U��]�u��e����ڋU����ց���  f;��]�U��f;�M����  f;�}B��������E�t�E��U��]�u��m�����ڋU������H�]�U�u�9E�tf�M�f�}� �w�U����� �� � u1�}��u(�}���E�uf�}����E�u	f�E� �G�f�E���E���E�f���rf�ىE�E�Ɂ�   ��� ���M�3��6f�E�f�E��E�E�E���E�f�}���f��Ɂ�   ��� ���M�E�E��E�U��M�f�
t2��M9E'f�" f�}� ��B����$ �B�B0�B ����jY9M~�M�u���j���?  f�E�[�E��}�M��e������E�����K�}�E�uڅ�}2�ށ��   ~(�E�}�M��m�������E������N���}�E�؋E@���Z�]��E���   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B�ҋ�tA�Eȍ0;։U�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K���K�K<5}�M��D�;9u	�0K;]�s�;]��E�sCf� �*؀��ˈX�D �E��M�_^3�[��x���À;0uK;�s�;ًE�s�f�  f�}� ��@���ʀ��� �P�0�@ �����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u�����   ^t   �3���t��   ��SVW�   t���t   ��t   ��t   ��   �   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#с�   ^[t��   t
;�u �  Ã�@�@�  Ã�SUVW��|$�\$3���tjZ��t����t����t���� t����t��   �ˋ��   #ǽ   �   t =   t=   t;�u��
����   #�t;�u��   ���   f�� t��   �t$(�L$$����#�#��;D$��   ���������D$�l$��|$�\$3���tjZ��t����t����t���� t����t��   �ˋ�#�t$=   t=   t;�u����   ���   #�t��   u��   ���   f�� t��   �T$�=�� ��  �����\$�D$3���yj^f� t��f� t��f� t��f� t��f� t��   �Ƚ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #Ã�@t-�  t��@u��   ���   ���   ��#|$$��#��;�u���   �"���P�D$,�k���Y�\$(�D$(3҄�yjZ�   ��t��f� t��f� t��f� t���   ��t��   ��#�t"��    t�� @  t;�u��   ����#Ã�@t-�  t��@u��   ���   ���   �L$��3���� t   �_^][���U���VW�u�M��B����E�u3�;�t�0;�u,�����WWWWW�    �kx�����}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP�`���M������   ���B����t�G�ǀ�-u�M���+u�G�E���I  ���@  ��$�7  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   ���3��u���N��t�˃�0�f��t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �\�]��]ى]��G댨����u�u>��t	�}�   �w	��u,9u�v'�.����E� "   t�M����E$�����ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^��U��3�9��P�u�u�uuh�-�P������]�U���SVW3�jSS�u�]��]���}���E�#�����U�tYjSS�u��}����#ʃ����tA�u�}+����   ;���   �   Sj�@ P�< ���E�u�"����    ����� _^[��h �  �u�  YY�E���|
;�r�����P�u��u��~�������t6�+��xӅ�wϋu��u��u��   YY�u�j �@ P�4 3��   �����8u�����    ����u��;�q|;�skS�u�u�u��|��#�����D����u�2_��YP�,!�����H��E�#���U�u)�6����    �>������D ��u�#u��������S�u��u��u�`|��#���������3������U��U������k�8S�]V�4������A%�   �E�A$���W� @  ��;�tP�� �  tB��   t&��   t��   u=�I���L$��⁀���'�I���L$��₀���a��I���L$�!��} u� �  ����% �  �_^[]ËD$V3�;�u�"���VVVVV�    ��s����jX^Ë(��3�^�3�PPjPjh   @h̶�!��5á�5���V�5� t���tP�֡�5���t���tP��^�U��QV�uV腒���E�F��Yu����� 	   �N ���  �;  �@t�w���� "   ��t�f ���   �N�����F�F�f �e� Sj���[�f��Fu,�ih���� ;�t�]h����@;�u�u�!�����YuV�ҷ��Yf�FW��   �F�>�H��N+�+˅��N~WP�u蛁�����E��N�� �F�?����M���t���t����k�8����������)�@ tSj j Q�pz��#����t-�F�]f��j�E�P�u���]f�]��#������E�9}�t�N ���  ���%��  _[^��U����  3ŉE��ESV3�9uW�E�N@  �0�p�p�F  ��X���}𥥥�����<�ыH�����Ή}���e� �������ˋ]���׍<;��0�P�Hr;�s�E�   3�9]�8t�r;�r��s3�C�ۉptA�H�H�U�3�;�r;�s3�F���Xt�@�M�H�e� �?�����<��P������Uމ�x�X��4;�U�r;�s�E�   �}� �0t�O3�;�r��s3�B�҉HtC�X�M�E�} �����3��&�H�����P�����������E���  �H�9ptջ �  �Xu0�0�x�E���  ������0�4?�H�����ʅˉp�Ht�f�M�f�H
�M�_^3�[�l������% �������̋D$�L$PQ�J�����������������̋D$P�J��Y����̋M������M���������M��� ������M���0������M���@������T$�B�J�3��k�����=h��̋M������M��������M��� �����M���0�����M���@�����T$�B�J�3��5k������g��̍M�h����E����   �e���M�P���ÍM��G����M��?����M��7����M��/����M��'����T$�B�J�3���j���(�g��h�#j}hD��E�P��3����ËT$�B�J�3��j�����Tg���������̋E����   �e���M����ËT$�B�J�3��`j�����g�������������̍�����e����M��}����M��u����M��m����M��e����M��]����M��U����������J����������?����������4����������)����� ��������� ���������@���������`����������p�����������������������������������������M��������0�������������������P���������p������������������T$�B�����3��8i������e�����̍M��h����E����   �e���M�P���ËT$�B�J�3���h�����e�����̍M�����E����   �e���M����ËT$�B�J�3��h����pe�����̍�t���������T$�B��P���3��h�����Ce���M������T$�B�J�3��hh���J�3��^h�����e���M������M������M�������d����w�����8����l�����(����a�����H����&����������������������������������H���������M�By���M������M������M��
�����t���������M�������M�������M��������,���鬟����d���顟��������閟��������鋟��������速���M�������t��������M������T$�B��(���3��;g������c���M��5���M��~�����������T$�B�����3��g���0�c���M��f5���M��n~����h����S���T$�B��L���3���f���l�c���M��M����l����"����M�������M�������M�������M�������M�������M�������M��
L���M�������M������T$�B��|���3��Pf�����c���M������M��|����T$�B�J�3��%f�����b���M��y~���T$�B�J�3��f���H�b���M��V~���T$�B�J�3���e���t�b����ȸ��� %����(�������������D�������������������w��������������������������д��铝���������������������������������������gP���M�������|����TP����@���������X����>P�������������������(P����`����m����������P��������G����������,���������A�����������O���M��.�����|�����O����8���������X����O����h����O����Զ�������������霜��������������@����������`����{O��������������������eO����`���������p����OO�������������� ����9O����\����~�����8����#O���������h�����P����O����<����R����������N��������<�����$�����N��������&����������N����|�������������N����,��������������N����L���������������N����l��������������sN��������������8�������������RN��������釆����ܸ���|����������a�����|����v���������N����$����`����������N����\����J����������M��������4����������M�������������������M��������������$����M�������������������M�������������������M����Ե��������������kM�������������4����UM�������������������?M����<���������t����)M��������n�����T����M����l����X�����4�����L����ĵ���B�����$�����L����L����,����������L����|���������D����L��������� ����������L����Զ���������d����L��������������h����yL����8��������������cL�������������H����ML�������������M��:L���������_����������$L���������i�����|����L����8����S�����X�����K��������=�����`�����K����Զ���'�����������w��������������M������������������������������������������������������������T$�B������3��X`���J�3��N`�����]�����������̋T$�B�J�3��)`������\�������h&jhD��E�P�+)����ËT$�B�J�3���_���H�\�������������̋M��`���T$�B�J�3���_���t�y\��������������̍M�鸂���T$�B�J�3��_�����I\��������������̋M��8`���T$�B�J�3��a_���$�\��������������̍M��X����T$�B�J�3��1_���P��[��������������̍M��(����T$�B�J�3��_���|�[��������������̋E���   �e���M����ÍM��/����E���   �e���M���I��ËT$�B�J�3��^�����W[���M�������M�������M��������d���������8���������(���������H����g����������\����������Q���������F�����H����;����M�o���M��[����M��S����M��K�����t����@����M��8����M��0����M��(�����,���������d��������������ו���������̕��������������M��������t���������M�������T$�B��(���3��|]�����4Z���M������M������M������T$�B�J�3��I]���0!�Z���M����T$�B�J�3��&]���\!��Y���M��z���M��r����M��j����M��H���M��
H���M��R����M���G���M��B����M���G���M�2���T$�B������3��\����!�pY����x��������M������T$�B��t���3��\���"�?Y���E�P��"��YÍ�8��������M������T$�B��t���3��K\���@"�Y���������~���������������������������{���������p����T����e�����L����
G�������������������D����T����9������������   ���������L�����F��Í�l���鼓�������鱓��������馓����<���������������������������   ���������4����oF��ÍM����������������$���������D����EF��������:F����l����/F�������������������i���������^��hp(h  hD�������P�$����Í�P����4���M�����hp(ho  hD���x���P��#����Í��������������������T����������$����������<���������\���������<���������|������hp(h�  hD�������P�Z#����Í�L����k����M��c�����<����X����T$�B������3���Y���J�3���Y���d"�V���EP�M�Q�#�����ËT$�B�J�3���Y����#�V�����̋EP�M�Q�������ËT$�B�J�3��Y���$�PV�����̋EP�M�Q�������ËT$�B�J�3��hY���8$� V�����̋EP�M�Q������ËT$�B�J�3��8Y���d$��U�����̋EP�M�Q�c�����ËT$�B�J�3��Y����$��U������hp(jhD��E�P�"����ËT$�B�J�3���X����$�U�������������̍M���{���T$�B�J�3��X����$�YU��������������̍M��{���T$�B�J�3��qX���%�)U��������������̍M��h{���T$�B�J�3��AX���P%��T��������������̍M��8{���T$�B�J�3��X����%��T��������������̍M��{���T$�B�J�3���W����%�T��������������̍M���z���T$�B�J�3��W��� &�iT��������������̍M��z���T$�B�J�3��W���,&�9T��������������̍�<��������T$�B��0���3��KW���X&�T��������̍M��x����E����   �e���M�`���ËT$�B�J�3��W����&��S�����̍����������������*���������o����������������������   ������������������Ë��������   ���������t��������Í������������t��������T$�B��H���3��`V���J�3��VV����&�S��h8*h�   hD��E�P�Z����ËT$�B�J�3��V���'��R������������̍M�H����M�@����T$�B��J�3���U���P'�R������̡�9�����9ËT$�B��J�3��U���|'�sR��������̡�9�����9ËT$�B�J�3��U����'�CR��������̋M������T$�B�J�3��aU����'�R��������������̋EP�M�Q������ËT$�B��J�3��(U��� (��Q�����̋E�P�w��YËT$�B��J�3���T���,(�Q�����������̋E�P�G��YËT$�B�J�3���T���X(�Q�����������̋M��X����M����   �*L���T$�B�J�3��T����(�KQ����������������̋M������T$�B��J�3��aT����(�Q��������������̋M������M���4�N���M���h����T$�B��J�3��T����(��P��������̋E�P�g��YËT$�B��J�3���S��� )�P�����������̋E�P�7��YËT$�B�J�3��S���L)�vP�����������̋E�P���YËT$�B�J�3��S���x)�FP�����������̋M��8����M���4�=M���M���h�����T$�B��J�3��KS����)�P��������̋E�P���YËT$�B��J�3��S����)��O�����������̋E�P�g��YËT$�B�J�3���R���*�O�����������̋EP�M�Q������ËT$�B��J�3��R���8*�pO�����̋M��xL���T$�B�J�3��R���d*�IO��������������̋M��8����M��������M��������M���,�wy���M����   �i���T$�B��J�3��2R����*��N���������������̋M�������M����m���M����b���M���,�y���M����   �)i���M����   ��l���T$�B�J�3���Q����*�|N���E�P���YËT$�B��J�3��Q���0+�VN�����������̋E�P����YËT$�B�J�3��nQ���\+�&N�����������̍M������T$�B��J�3��AQ����+��M��������������̋E����   �e���M�X���ËT$�B�J�3�� Q����+�M�������������̍M��(����T$�B��J�3���P����+�M��������������̍M�������T$�B��J�3��P���,�YM��������������̍�����������T$������������3��hP���8,� M�����̍�0���������`������������������T$������������3��"P���t,��L���������������̍M��8���E�P���YÍM��Ճ���T$��L�����H���3���O����,�L�����̍M������T$�BȋJ�3��O����,�iL��������������̍M�������T$�B��J�3��O���-�9L��������������̍M������M������T$�B��J�3��IO���<-�L������̋E�P���YËE�P���YËT$�BЋJ�3��O���p-��K����������������̋E�P�W��YËT$�B�J�3���N����-�K�����������̋E�P�'��YËT$�B��J�3��N����-�fK�����������̋M������T$�B�J�3��N����-�9K��������������̋M�������T$�B��J�3��QN��� .�	K��������������̋M������T$�B��J�3��!N���L.��J��������������̍M��x����M��p����T$�B��J�3���M����.�J������̍M��H����T$�B��J�3���M����.�yJ��������������̍�X���������M�������h��������T$����������3��uM����.�-J��̍�8��������T$����������3��HM���/� J�����̍M��x����T$�B�J�3��!M���@/��I��������������̍M�H����T$�B�J�3���L���l/�I��������������̍M������T$�B�J�3���L����/�yI��������������̍�\����E���T$��\�����X���3��L����/�@I�����̍�P��������T$����������3��XL����/�I�����̍�0��������T$����������3��(L���0��H�����̋EP�w��YËT$�B�J�3���K���H0�H�����������̍������%����T$������������3���K���t0�H�����̍M�������T$�B�J�3��K����0�YH��������������̍M�������T$�B�J�3��qK����0�)H��������������̍�(��������T$����������3��8K����0��G�����̍M��h����T$�B��J�3��K���$1��G��������������̍�`����5���������Z�����H����~���T$������������3���J���`1�zG���������������̍������%b����H����������8���������T$������������3��rJ����1�*G���������������̍�x���������������	����d����a���������t����T$��L�����H���3��J����1��F����̍������E����T$������������3���I���2�F�����̍������U���������:���������?���������$���T$��L�����H���3��I���P2�OF����̋M��X���T$�B�J�3��qI���|2�)F��������������̍�����������8�����`����`���������@����t����T$����������3��I����2��E����̍�8��������T$��<�����8���3���H�����J�3���H����2�E��������̋M��h����T$�B܋J�3��H���3�iE��������������̋M���0������T$�B�J�3��~H���D3�6E�����������̍M�����T$�B��J�3��QH���p3�	E���������������h@jj�E�P�s��ËT$��L�����H���3��H����3��D�������������̍M��8����T$�B��J�3���G����3�D��������������̋E����   �e���M�����ËT$�B��J�3��G����3�XD�������������̋E�P����YËT$�B��J�3��nG��� 4�&D�����������̋E�P���YËT$�B�J�3��>G���L4��C�����������̋E�P���YËT$�B��J�3��G���x4��C�����������̋E�P�W��YËT$�B�J�3���F����4�C�����������̋E�P�'��YËT$�B��J�3��F����4�fC�����������̋E�P����YËT$�B�J�3��~F����4�6C�����������̋M������T$�B��J�3��QF���(5�	C��������������̋E�P���YËT$�B��J�3��F���T5��B�����������̋E�P�g��YËT$�B��J�3���E����5�B�����������̋EP�7��YËT$�B�J�3��E����5�vB�����������̋EP�M�Q�������ËT$�B��J�3��E����5�@B�����̋M����Ud���T$�B�J�3��^E���6�B�����������̋Eă��   �e���M�x���ÍM��/K���T$�B��J�3��E���86��A�����̍�8���镽���T$��4�����0���3���D�����J�3���D���d6�A��������̋M��h����M����   �*���T$�B�J�3��D����6�[A����������������̋M�����[���M����:b���M���$�ob���M���4�b���T$�B��J�3��MD����6�A����������̍M��x����T$�BȋJ�3��!D���7��@��������������̍M��H����T$�BȋJ�3���C���47�@��������������̋E�P�7
��YËT$�B��J�3��C���`7�v@�����������̋E�P�
��YËT$�B�J�3��C����7�F@�����������̋E�P��	��YËT$�B�J�3��^C����7�@�����������̍����酾���M��}����T$����������3�� C����7��?�������������̍M��8���T$�BȋJ�3���B���8�?��������������̍�����������p����
����T$������������3��B���L8�e?����������̋M��#���M����͆���M�����a���M���(������M���8�����M����   �����M����   �����M���   �2Y��h@jj�E�  P�m���h@jj�E�@  P�m��ËM���d  �db���M���  �v_���M���   �^���M���8  �ʚ���T$�B�J�3���A���p8�{>����������������̋M��"���M����݅���M����a���M���(�����M���8������M����   �.����M����   �����M���   �BX��h@jj�E�  P�l���h@jj�E�@  P�l��ËM���d  �ta���M���  �^���M���   �]���M���8  �ڙ���T$�B�J�3���@���9�=����������������̋E�P���YËT$��L�����H���3��@����9�P=�����̋E�P����YËT$�B��J�3��n@����9�&=�����������̋E�P���YËT$�B�J�3��>@����9��<�����������̋M��(!���M����]����M����_���M���(釄���M���8�|����M����   鮄���M����   � ����M���   ��V��h@jj�E�  P�=k���h@jj�E�@  P�%k��ËM���d  ��_���M���  �]���M���   �(\���M���8  �Z����T$�B��J�3��S?���:�<����������������̋E�P���YËT$�B�J�3��?����:��;�����������̋M�� ���M����=����M����b^���M���(�g����M���8�\����M����   鎃���M����   � ����M���   �U��h@jj�E�  P�j���h@jj�E�@  P�j��ËM���d  ��^���M���  ��[���M���   �[���M���8  �:����T$�B�J�3��3>����:��:����������������̍M�x����T$�B��J�3��>���x;�:��������������̋M������M����   �����T$�B�J�3���=����;�{:����������������̋M�����T$�B��J�3��=����;�I:��������������̍M�鸸���T$�B��J�3��a=���<�:��������������̋M������M����   �����T$�B�J�3��#=���8<��9����������������̋M�騚���M����   �Z����T$�B�J�3���<���l<�9����������������̋E�P�'��YËT$�B��J�3��<����<�f9�����������̋E�P����YËT$�B�J�3��~<����<�69�����������̋E�P����YËT$�B��J�3��N<����<�9�����������̋E�P���YËT$�B�J�3��<���=��8�����������̋E�P�g��YËT$�B�J�3���;���H=�8�����������̍M��8����T$�B�J�3���;���t=�y8��������������̋M�����M���������M���(������M���,������M���0������M���4������M���@馶���M���p�@���M����   �����M����   �_����T$�B��J�3��(;����=��7�����̋M�����M����]����M���(�b����M���,�W����M���0�L����M���4�A����M���@�����M���p�@���M����   �����T$�B��J�3��:���>�^7���̍M�������T$�B�J�3��:����>�97��������������̍M������M������T$�B܋J�3��I:����>�7������̋M��ؗ���M����   �����M����   �����T$�B��J�3��:����>�6��̋M�阗���M����   �z����M����   �ܵ���T$�B��J�3���9���,?�}6��̋E�P� ��YËT$�B��J�3��9���X?�V6�����������̋E�P�����YËT$�B�J�3��n9����?�&6�����������̋E�P����YËT$�B��J�3��>9����?��5�����������̋M�������M���4��2���T$�B�J�3��9����?�5���̋EP�W���YËEP�L���YËT$�B�J�3���8���@�5����������������̋E�P����YËT$�B�J�3��8���D@�V5�����������̍M��ȳ���M�������M�鸳���T$�B��J�3��a8����@�5��������������̍�@���酳���T$������������3��(8����@��4�����̋M������M����M����M���8�B����M����   �4����T$�B�J�3���7����@�4����������̋M�����M���������M���8�����M����   �����T$�B��J�3��7���4A�E4����������̍M�鸲���T$�B��J�3��a7���`A�4��������������̍M�鈲���T$�B��J�3��17����A��3��������������̍�0����U����������J����T$��L�����H���3���6����A�3����������̍M������M�������d��������T$��h�����d���3��6����A�`3�����̋EЃ��   �e���M��ȱ��ËEЃ��   �e���M鯱��ËT$�BԋJ�3��W6���0B�3����̍M������T$�B��J�3��16���\B��2��������������̋�����P�t���YËT$��L�����H���3���5����B�2��̍M��(����T$�B��J�3���5����B�2��������������̍������%��������������T$������������3��5����B�E2����������̍�,���鵰���� ���P�����YÍ�,���霰���� ���P����YË� ���P����YËT$����������3��#5���C��1����������������̋EP�g���YËT$�B�J�3���4���`C�1�����������̋EP�M�Q������ËT$�B��J�3��4����C�p1�����̋EP�M�Q������ËT$�B��J�3��4����C�@1�����̋EP�M�Q賯����ËT$�B��J�3��X4����C�1�����̋EP�M�Q胯����ËT$�B��J�3��(4���D��0�����̋M�������M����M����M���8�B����M����   �4����T$�B��J�3���3���TD�0����������̍�H��������M��������(���������8���������$���P�����YËT$����������3��|3���xD�40���������̍�����饮����@���隮����p���鏮�������鄮���� ����y�����0����n����� ����c���������P�w���YË�����P�i���YË�����P�[���YË�����P�M���YËT$������������3���2����D�/�����������̋M��X����T$�B�J�3��2���HE�Y/��������������̋M��(����T$�B��J�3��q2���tE�)/��������������̋E�P����YËT$�B��J�3��>2����E��.�����������̋E�P����YËT$�B�J�3��2����E��.�����������̋E�P�W���YËT$�B��J�3���1����E�.�����������̋E�P�'���YËT$�B�J�3��1���$F�f.�����������̍������K��������������`����7��������P�����YËT$������������3��T1���hF�.���EP����YËEP����YËEP����YËT$�B�J�3��1����F��-�����̍M��H�����|����=����T$��|�����x���3���0����F�-�������������̍�T����������@����������0���������p��������T$������������3��0���G�?-����̍M�鸫���T$�BċJ�3��a0���HG�-��������������̍M�鈫���T$�B��J�3��10���tG��,��������������̋E����   �e���M��H���ËE����   �e���M��/���ËT$��|�����x���3���/����G�,��������������̍M�����T$�B�J�3��/����G�Y,��������������̍M��Ȫ���M�������T$�B��J�3��i/���H�!,������̍�h���镪����X���銪���T$����������3��-/���<H��+����������̍M��X����T$�B��J�3��/���hH�+��������������̍M��(����T$��L�����H���3���.����H�+��������̍�`���������M������T$��\�����X���3��.����H�H+�������������̍�`���鵩���M�魩���T$��T�����P���3��P.����H�+�������������̍�0����u����T$������������3��.���(I��*�����̋M������T$�B��J�3���-���TI�*��������������̋M��h����T$�B��J�3���-����I�y*��������������̋M��8����M���p�����M����   �Ϩ���T$�B�J�3��x-����I�0*�����̋M�������M���p魶���T$�B��J�3��F-����I��)���̋M��8���M����mD���T$�B�J�3��-���$J��)���̋M�����M����=D���T$�B��J�3���,���XJ�)���̋M������M����D���M���H�����T$�B�J�3��,����J�c)��������̋M��X����M�����C���M���H�§��h@jj�E���xP��W��ËT$�B��J�3��U,����J�)��̍�����酧���������z����T$������������3��,���K��(����������̍M��H����T$�B��J�3���+���8K�(��������������̍����������������
�������������������������h@jj������P�!W��Í������Ӧ���T$��L�����H���3��v+���\K�.(���̍�8���饦����p���隦���T$����������3��=+����K��'����������̍M��X����T$�BԋJ�3��+����K��'��������������̍M��(����T$�BԋJ�3���*���L�'��������������̍M�������T$�BԋJ�3��*���DL�i'��������������̍M������T$�B��J�3��*���pL�9'��������������̍M�������T$�BȋJ�3��Q*����L�	'��������������̍M��x����M��p����M��h����M��`����T$�B��J�3��	*����L��&������̍M��8����M��0����M��(����M�� ����T$�B��J�3���)���$M�&������̋EP�M�Q������ËT$�B�J�3��)���PM�P&�����̋E�P�����YËT$�B�J�3��n)���|M�&&�����������̋E�P����YËT$�B��J�3��>)����M��%�����������̋E�P����YËT$�B��J�3��)����M��%�����������̋E�P�W���YËT$�B�J�3���(��� N�%�����������̋E�P�'���YËT$�B��J�3��(���,N�f%�����������̋E�P�����YËT$�B�J�3��~(���XN�6%�����������̍M�騣���T$�B��J�3��Q(����N�	%��������������̋E�P����YËT$�B��J�3��(����N��$�����������̋E�P�g���YËT$�B�J�3���'����N�$�����������̋E�P�7���YËT$�B��J�3��'���O�v$�����������̋E�P����YËT$�B�J�3��'���4O�F$�����������̍�����鵢��������骢����x���韢��������锢��������鉢����x����~���������s����������h����������]���������R����M��J����M��B����T$������������3���&���XO�#��̋E�P�M�Q������ËT$�B�J�3��&����O�p#�����̋E�P�M�Q������ËT$�B�J�3��&���P�@#�����̋E�P�M�Q賡����ËT$�B�J�3��X&���<P�#�����̋E�P�M�Q胡����ËT$�B�J�3��(&���hP��"�����̍M��X����T$�B܋J�3��&����P�"��������������̋M������M�������M��� ����M���0����M���@�z���M���P�z���M���`�z���M���p�z���M����   �z���M����   鿠���T$�B��J�3��h%����P� "�����̋M��X���M��������M��� �����M���0�����M���@�z���M���P�!z���M���`�&z���M���p�+z���M����   �-z���M����   �/����T$�B��J�3���$���,Q�!�����̍M������M�� ����T$�BЋJ�3��$����Q�a!������̍�T����՟����D����ʟ����d���鿟����d���鴟���T$��@�����<���3��W$����Q�!����̍�D���酟����4����z�����d����o�����T����d����T$��8�����4���3��$���8R� ����̍M�8����M�0����������%����������������������������������T$������������3��#���\R�_ ����̍M��؞���M��О���T$�BԋJ�3��y#����R�1 ������̍M������T$�BԋJ�3��Q#����R�	 ��������������̍M��h����T$�BЋJ�3��!#��� S����������������̍M��8����T$�BЋJ�3���"���TS���������������̍M������T$�BЋJ�3���"����S�y��������������̍M�������T$�B̋J�3��"����S�I��������������̍M��(?���T$�BȋJ�3��a"����S���������������̍M�鈝���M�逝���M��x����M��p����T$�B��J�3��"���T��������̋E�P�g���YËT$�B��J�3���!���HT������������̋E�P�7���YËT$�B�J�3��!���tT�v�����������̋E�P����YËT$�B��J�3��!����T�F�����������̋M��x���M�������M��� ����M���0����M���@�<v���M���P�Av���M���`�Fv���M���p�Kv���M����   �Mv���M����   �O����T$�B�J�3��� ����T������̍M��(����T$�B��J�3��� ���@U���������������̍M�������T$�B��J�3�� ���lU�Y��������������̍�D��������T$����������3��h ����U� �����̋EP����YËT$�B��J�3��> ����U�������������̋M��(���T$�B��J�3�� ����U����������������̋E�P�W���YËT$�B��J�3������V������������̋E�P�'���YËT$�B�J�3�����HV�f�����������̋M��h{���T$�B��J�3�����tV�9��������������̋M��8{���T$�B��J�3��Q����V�	��������������̋M�����F���T$�B��J�3������V�������������̋M��h����T$�B�J�3�������V���������������̋EP�M�Q������ËT$�B��J�3�����$W�p�����̋EP�M�Q������ËT$�B��J�3�����PW�@�����̋EP�M�Q賙����ËT$�B��J�3��X���|W������̋EP�M�Q胙����ËT$�B��J�3��(����W�������̋EP�M�Q�S�����ËT$�B��J�3�������W������̋EP�M�Q�#�����ËT$�B��J�3������ X������̋EP�M�Q������ËT$�B��J�3�����,X�P�����̋EP�M�Q�Ø����ËT$�B��J�3��h���XX� �����̋EP�M�Q蓘����ËT$�B��J�3��8����X�������̋EP�M�Q�c�����ËT$�B��J�3������X�������̋EP�M�Q�3�����ËT$�B��J�3�������X������̍M��(����M�� ����M������T$�B܋J�3�����Y�Y��������������̍M�������T$�B��J�3��q�����J�3��d���DY����M���D�%����M���T�����M���d�����M���t�����M����   ������M����   ������T$�B��J�3�����hY���������������̍�D����E����T$��@�����<���3��������J�3������Y�s��������̍M������T$�B��J�3������Y�I��������������̍M�������T$�B��J�3��a�����J�3��T���Z����M������T$�B��J�3��1���HZ����������������̍M������T$�B��J�3�����tZ���������������̍M��X����T$�B��J�3�������Z���������������̍�8����E����T$��4�����0���3�������J�3������Z�C��������̍M���(���T$�B��J�3��a�����J�3��T����Z����M��H����T$�BЋJ�3��1�����J�3��$���$[��������������T$������������3��������J�3������P[���������̍�(�������T$��$����� ���3�������J�3�����|[�c��������̍�(����%����T$��$����� ���3��x�����J�3��k����[�#��������̋M��(u���M����@���T$�B�J�3��6����[�����̍M��h0���T$�B܋J�3�����x\����������������̍M������T$�B��J�3��������J�3�������\�����X����E����T$��T�����P���3�������J�3������\�S��������̋M����U����M�����0���M����   �y���M����  �����M����  �@���M����  �b���M����  �����M����  ����M����  ����M���  �J���M���  �L���M���(  �4���M���8  �@���M���H  �B���M���X  �T4���M���h  �����M���x  �4���M����  �j����M����  �\����M����  �N����M����  �@����M����  颒���T$�B�J�3��K����\���������̋M��������M����/���M����   ��w���M����  �>����M����  �����M����  ����M����  �t���M����  �6���M����  �����M���  �����M���  �����M���(  ��2���M���8  �����M���H  �����M���X  �3���M���h  �f����M���x  �H3���M����  �����M����  �����M����  ������M����  �����M����  �R����T$�B��J�3�������]���������̍M������T$��|�����x���3��������J�3������^�v�����������̍���������������:����������
���T$������������3��r�����J�3��e����^���̋M���D�%����M���T�����M���d�����M���t�����M����   ������M����   ������M����   ������T$�B��J�3������_�����������������̍�@��������T$��H�����D���3�����h_�p�����̍M������T$�B��J�3�������J�3������_�<���������e���������P�����YÍ������L���������P����YÍ������3���������P����YÍ���������������P�~���YÍ���������������P�e���YÍ����������������P�L���YÍ������������8����t;������������������P����YÍ���������������������8����:;���������%���T$������������3��r�����J�3��e����_���̋M��X����M��������T$�B��J�3��6����`�����̋M��(����T$�B��J�3������`����������������̋E�P�W���YËT$�B��J�3�������`������������̋E�P�'���YËT$�B�J�3�����a�f�����������̍� ���������@����ʍ���������������P���鴍���T$����������3��W���4a�����̋M������M��������T$�B��J�3��&����a�����̋M��ب���M����m����T$�B��J�3�������a����̋M�騨���M����=����M����   �����T$�B��J�3����� b�p�����̋M��h����M���������T$�B��J�3�����4b�>���̍M��+���T$�B؋J�3��a���`b���������������̍M�����T$�B��J�3��1����b����������������̋E�P�w���YËT$�B��J�3�������b������������̋E�P�G���YËT$�B�J�3�������b������������̋E�P����YËT$�B��J�3�����c�V�����������̋E�P�����YËT$�B�J�3��n���<c�&�����������̋M�����)���T$�B��J�3��>���hc�������������̋M������M����}����M��� �r����M���d釺���M���t�l����T$�B�J�3�������c���̋M�阦���M����-����M��� �"����M���d�7����T$�B��J�3������c�X�������������̋E�P�����YËT$�B��J�3��n���$d�&�����������̋E�P����YËT$�B�J�3��>���Pd�������������̋M������T$�B��J�3�����|d����������������̍M��X����T$��L�����H���3�������d���������̋M�����M�����M�����4���T$�B��J�3������d�V�����������̋M������T$�B��J�3��q���e�)��������������̋E�P����YËT$�B��J�3��>���<e��
�����������̋E�P����YËT$�B�J�3�����he��
�����������̍�@����5����T$����������3�������e�
�����̍�@��������T$����������3������e�`
�����̍M�������T$�B�J�3������e�9
��������������̋M���(������T$�B��J�3��N���f�
�����������̋M���(�����T$�B��J�3�����Df��	�����������̋M��H����T$�B��J�3������pf�	��������������̋M������T$�B��J�3�������f�y	��������������̍M������T$�B��J�3�������J�3������f�<	���M�鸇���T$��`�����\���3��[�����J�3��N����f�	�����������̋M���x�����M���|�����M����   �|����T$�B��J�3�����0g���̋EP�M�Q�3�����ËT$�B��J�3������\g������̋M��� �%����M���$�����M���(�����M���,�����M���0������M���4������M���8������M���<������M���@������M���D������T$�B��J�3��K����g���������̋M���d�����T$�B��J�3������g�������������̋M��H����M����   �Z����T$�B��J�3���
���0h�����������������̋M������M����   �����T$�B�J�3��
���dh�[����������������̋M�������T$�B��J�3��q
����h�)��������������̋M���8�����T$�B�J�3��>
����h�������������̋M���x�����M���|�z����M����   �l����M����   �^����T$�B��J�3���	��� i�����̋EP�M�Q������ËT$�B��J�3��	���,i�p�����̋M��(����M���(  ��X���M���X  ������M����  ��&���M����  �@���M����  ��#���M���   �$����T$�B�J�3��=	���Pi������������̋M������M���(  �zX���M���X  �l����M����  �^&���M����  �����M����  �r#���T$�B��J�3�������i���������̋M�������E�P�M�Q������ËT$�B�J�3�����j�H�������������̍�T����E���T$��P�����L���3��X���<j������̋E�P�M�Q胃����ËT$�B�J�3��(���hj�������̋M��x����M��� �4���M����   �?���M����   �1���M���  �#����M����  �����M����  �����M���P  �����M����  �^���M����  �-f���M����  �f���M���(  �����M����  ��a���T$�B�J�3��\����j����������̋M������M��� �=3���M����   �o���M����   �a���M���  �S����M����  �E����M����  �7����M���P  ����M����  �]���M����  �]e���M����  �Oe���M���(  ����T$�B��J�3�����k�R�������̍������uZ���T$������������3��h�����J�3��[����k���������̍������5Z���� ����
���������Z���T$������������3�������J�3������k���̋E����   �e���M�(���ËT$�B�J�3������l��������������̍M�����T$��J�3�����8l�Z���������������̋M����U����T$�B��J�3��n���dl�&�����������̋M���b���M����   銀���T$�B�J�3��3����l������������������̋M��b���T$�B��J�3������l���������������̋EP�M�Q�#�����ËT$�B��J�3�������l������̋EP�M�Q������ËT$�B��J�3�����m�P�����̋E�P�����YËT$�B��J�3��n���Hm�&�����������̋E�P����YËT$�B��J�3��>���tm�� �����������̋E�P�M�Q�c����ËT$�B�J�3������m�� �����̋M��� 酛���T$�B�J�3�������m� �����������̋M��� �U����M����@  �����T$�B�J�3����� n�X �������������̍M���~���E�P�����YËT$�B��J�3��f���4n� ���̍M��~���E�P����YËT$�B��J�3��6���hn������̋M��Ȱ���T$�B�J�3������n�����������������̋M�阰���T$�B�J�3�������n����������������̋E�P�M�Q�~����ËT$�B�J�3������n�`������̋E�P�M�Q��}����ËT$�B�J�3��x���o�0������̍M��8����T$�B̋J�3��Q���Do�	���������������̍M������EP����YËT$�B؋J�3�����xo������̍M��ء���M��С���M��ȡ���M�������M�鸡���M�鰡���T$�B��J�3�������o��������̋M��x����M��������M��� �����M���d�����T$�B�J�3�����p�8��������������̍� ���������P���P����YËT$��L�����H���3��:�����J�3��-���Dp�������������̍M������EP�o���YËEP�d���YËEP�Y���YËEP�N���YËT$�B��J�3��� ���hp����̍�0����%�����8���P����YÍ�h�����{����8���P� ���YÍ�h�����{����@����x����8���P�����YÍ�h����{����@����T����8���P����YÍ�h����{����@����0����8���P����YÍ�h����g{����@�������T$��,�����(���3���������J�3��������p�����������������̍M��{���E�P�/���YËT$��P�����L���3��������J�3������`q�[�����������������̍M���z���E�P�����YËE�P�����YËT$��L�����H���3��U�����q����̍M��x����M��z���T$�B��J�3��)�����q���������̍M��H����M��Pz���T$�B��J�3�������r��������̋EP�G���YËT$�B��J�3�������8r�������������̋EP����YËT$�B��J�3������dr�V������������̋E�P�����YËT$�B̋J�3��n�����r�&������������̋E�P����YËT$�BċJ�3��>�����r��������������̋E�P����YËT$�B؋J�3�������r��������������̋�x���P�T���YÍ�d����'y����d����y���M��y���T$��P�����L���3������,s�o�����̋E�P�M�Q��x����ËT$�B�J�3������Xs�@������̍�8����e������������������������T$����������3��B������J�3��5�����s�����̍���������T$������������3��������J�3��������s����������̍M�鸜���T$�B�J�3��������s����������������̍�X����5�����4���P�	���YËT$��$����� ���3��������J�3��}���� t�5�����������̍�����՘��������jl����P���������P����T����P��������P�������� ����C���T$����������3��������J�3�������Dt��������̍M鸛���T$�B��J�3��������t����������������̋E�P����YËT$�B�J�3�������t�V������������̍M������T$�B̋J�3��q���� u�)���������������̋M����%����M��������M��������M��������M���������M��� �����M���$�����M���(�ؚ���M���,�͚���T$�B��J�3�������$u�����̍M�騚���M頚���M�阚���M鐚���M�鈚���M�通���T$�B�J�3�������u�Q�������̍M��X����M�P����M��H����M�@����M��8����M��0����T$�B�J�3��I�����u��������̍M�����T$�B��J�3��!����@v�����������������̍M��ؙ���T$�B��J�3�������lv����������������̋M���饙���M���隙���M���鏙���M���鄙���M����y����M��� �n����M���$�c����M���(�X����M���,�M����M���0�B����T$�B��J�3��[�����v����������̍M��t���T$�B��J�3��1����w�����������������̋E����   �e���M�Ht��ËT$�B�J�3�������8w���������������̍M��t���M��t���T$�B��J�3������lw�q�������̍M������T$�BȋJ�3�������w�I���������������̍M������T$�BȋJ�3��a�����w����������������̍M�鸔���T$�BȋJ�3��1�����w�����������������̍������Us���T$������������3�������x�������̍������%s���������s����x����s����8����s����H�����r���������r����x�����r���T$��L�����H���3������@x�>����̍�0����r���T$����������3��X�����x�������̋E����   �e���M��xr��ËT$�B��J�3�� �����x����������������̋M��x����T$�B�J�3��������x����������������̋M��H����M����=����T$�B��J�3������0y�n����̋E�P����YËE�P�����YÍM���q���M���q���T$�B��J�3��s����ty�+�����������������̋E�P跼��YËT$�B��J�3��>�����y��������������̋E�P臼��YËT$�B�J�3�������y��������������̍�p����5q���M��]�����`����b����P����G����T$����������3������z�r��������̋M������M���������T$�B�J�3������Dz�>����̋M��ش���T$�B��J�3��a����pz����������������̋M�騴���M���靴���T$�B��J�3��&�����z������̋M��x����M����m����M����b����T$�B��J�3��������z����������̋M��h���M���T�	���M���p�����M����   �t���T$�B��J�3������${�U�����������̋M������M����ݳ���T$�B��J�3��f����X{�����̋M������M���T����M���p�����M����   ��
���T$�B��J�3�������{�������������̍M��Ho���T$�B��J�3��������{����������������̋E����   �e���M�o��ËT$�B�J�3�������{�h��������������̍M���n���T$�B��J�3������ |�9���������������̋E�P�ǹ��YÍM��͏���T$��L�����H���3��@����T|����������������̋E�P臹��YËT$�B��J�3�������|��������������̍M��8n���M��0n���M��(n���M��P����T$�B��J�3��������|��������̍M��(����T$�BċJ�3�������|�Y���������������̍M���-���T$�B܋J�3��q����}�)���������������̍M��m���M��m���T$�B��J�3��9����P}���������̍M��hm���T$��L�����H���3������|}�����������̍M��h����M��`����T$�B��J�3��������}��������̍M��m���T$�B��J�3�������}�i���������������̍M���l���M�� ����M��������`���������P���P�ѷ��YË�T���P�÷��YËT$��L�����H���3��D���� ~������������ul���M��ml���M��el���T$������������3������l~��������̍������5l���T$������������3��������~�������̋E�P�'���YËT$�B��J�3�������~�f������������̋E�P�����YËT$�B�J�3��~�����~�6������������̋E�P�Ƕ��YËT$�B��J�3��N�����������������̋M������T$�B��J�3��!����H�����������������̋M������T$�B��J�3�������t����������������̍�x����k���M��k����H����k���T$��<�����8���3��������]���̋E����   �e���M��j��ËT$�B�J�3��p������(��������������̍M��j���T$��L�����H���3��;����������������̍������ej���M��]j���M��Uj���T$������������3�������D��������̋M���0���T$�B��J�3�������p�����������������̍M���i���M���i���M���i���T$�B��J�3���������I���������������̍M��i���T$�B�J�3��a����؀����������������̋E�P觴��YËT$�B��J�3��.�������������������̋E�P�w���YËT$�B�J�3�������0��������������̋M��ȹ���M���(�i���T$�B��J�3�������d��~����̋M�阹���M���(��h���T$�B��J�3���������N����̍M�������M��������|�����x���T$��l�����h���3��X����ԁ�������̋E�P觳��YËT$�B��J�3��.���� ���������������̍M��Xh���T$�B��J�3������,�����������������̋M��ȸ���M؃��h���M؃�@�h���M؃�P�h���T$�B��J�3������p��h��������������̋M��x.���T$�B��J�3���������9���������������̍�����������p������������������T$������������3��2����؂������������������̍�����镸����p���骫�������韚���T$������������3�������������������������̍�p����E�����`�����f����(����O�����`���P����YËT$����������3������X��<�����@����f����0����f����`����f���T$����������3��B������������������������̍�0����ef����@����Zf���M��Rf���T$����������3�������Ѓ����̍������e�����p����z���������o����T$������������3��������j����������������̍�t�����e���T$��D�����@���3��x����8��0������̋E����   �e���M�e��ËT$�B�J�3��@����d�����������������̍M��he���T$��L�����H���3�������������������̋E�P�W���YËT$�B��J�3����������������������̋E�P�'���YËT$�B�J�3��������f������������̋M��x����M�����d���M���@��d���M���P�d���M���h�d���T$�B��J�3��U���������̍�����鵅��������骅����(����Ϩ��������tt���T$������������3������x�������̍�0����5d���� ����*d����@����d����P����d����`����	d�������P����YË����P����YËT$������������3���������H��������������̍�0����c����`����c���� ����c��������Ķ����@��������T$����������3��,������������������̍�8����Uc���T$����������3�������L��������̍�d����U����������z�����(����o����T$��L�����H���3���������j����������������̍M���b���M���b���T$�B��J�3��y�������1�������̍M��b���M��Ѓ���T$��L�����H���3��C�������������������������̍M��hb���M��`b���T$�B��J�3��	����$����������̍M��8b���M��0b���T$�B��J�3�������X���������̍M��b���M�� b����`�����a���M���a���M���a���M���a���M���a���M���a����p�����a���M��a���M��a����P����a���T$��L�����H���3��J����|����������̋M�騕���T$�B�J�3��!����������������������̋M��x����M��������T$�B�J�3�������<������̋M��H����M����}����M����B����T$�B�J�3������x��c���������̍M���`���T$�B��J�3���������9���������������̋E����   �e���M�`��ËT$�B�J�3��@����Ј����������������̍M��h`���M��``���T$�B��J�3��	��������������̍�(����5`���������*`���������`���������`���T$������������3������H��o�����̍������_����������_����@�����_���������_���T$������������3��g������������̍M��_���M��_���T$��L�����H���3��3�������������������������̍M��X_���T$��L�����H���3������������������̋E�P�G���YËT$�B��J�3���������������������̋E�P����YËT$�B�J�3������D��V������������̍M���^���M���^���M��^���M��^���M��8�����p���������T$��L�����H���3��@����h�����������������̍M��h^���M��`^���M�鈱����p��������T$��L�����H���3�������܊���������������̍M��^����8����^����h����^���M�銮���M��2�����(�����]����x�����]����X�����]����H�����]���T$����������3��i���� ��!�������̍M��]���M��]���M��]����\���������8���������l���������H���������0���P�p���YË�0���P�b���YËT$����������3�������l�������������������̍M�]���M�� ]���M���\���M���\���T$�B��J�3���������Q�������̍M������M��P����M��\���T$��L�����H���3��[����4�����������̍M��\����x����}\����P����r\���T$��L�����H���3������p������̋E�P�g���YËT$�B�J�3����������������������̋M��w���T$�B�J�3�������Ȍ�y���������������̍M�����T$�B��J�3��������I���������������̋M������T$�B�J�3��a���� �����������������̋M�騟���T$�B��J�3��1����L������������������̋M��x����T$�B��J�3������x�����������������̋E�P�G���YËT$�B��J�3����������������������̋E�P����YËT$�B�J�3������Ѝ�V������������̍�L����eD���T$��L�����H���3��h������J�3��[����������������̋E�P觥��YËT$�B��J�3��.����(���������������̋E�P�w���YËT$�B�J�3�������T��������������̋M��<���M����   �����T$�B�J�3����������{�����������������̋M��H<���T$�B��J�3���������I���������������̋E�P�פ��YËT$�B��J�3��^�������������������̋E�P觤��YËT$�B�J�3��.�������������������̍M��XY���M��PY���T$�B��J�3�������@���������̍M��X����T$�B�J�3�������l�����������������̍M������T$�B��J�3���������Y���������������̋M��(;���T$�B�J�3��q����ď�)���������������̍�@����X���T$������������3��8��������������̋M��(����M���$�}����T$�B��J�3������$������̋M�������M���$�M����T$�B��J�3�������X������̋M��h:���T$�B��J�3���������i���������������̋M��8:���M����   �����T$�B�J�3��s�������+�����������������̋M���9���T$�B�J�3��A����������������������̋M���9���T$�B�J�3������������������������̋E�P�W���YËT$�B��J�3�������<��������������̋E�P�'���YËT$�B�J�3������h��f������������̍�������V���T$����������3��x�������0������̍������V���T$������������3��H������� ������̋E�P藡��YËT$�B��J�3���������������������̋E�P�g���YËT$�B�J�3���������������������̍�h����V���T$��L�����H���3������D��p������̍M���U���T$��L�����H���3������p��C���������̍�����U���T$����������3��X�������������̋E�P觠��YËT$�B��J�3��.����Ȓ��������������̋E�P�w���YËT$�B�J�3����������������������̋EP�G���YËT$�B�J�3������� ��������������̋E�P����YËT$�B��J�3������L��V������������̋E�P����YËT$�B�J�3��n����x��&������������̋E�P跟��YËT$�B��J�3��>��������������������̋E�P臟��YËT$�B�J�3������Г��������������̋M�������M����-T���M����   ������M����   顅���T$�B��J�3��������r��������̍M������T$�B��J�3������@��I���������������̍M��S����X����ݦ���T$��L�����H���3��P����t����������������̍M�騦���T$�B��J�3��!�����������������������̍M��HS����X����m����T$��L�����H���3�������Ԕ���������������̍M��8����T$�B��J�3������ ��i���������������̍�(�����R����X����*����T$��$����� ���3��m����4��%�����������̍�\���������T$��\�����X���3��8����`���������̍M��hR����h���鍥���T$��L�����H���3�� ���������������������̍M��X����T$�B��J�3�������������������������̍M��(����T$�BЋJ�3��������Y���������������̍M���Q����h��������T$��L�����H���3��`���� ����������������̍M�鸤���T$�B��J�3��1����L������������������̋M������M����MQ���M����   ������M����   ������T$�B�J�3������������������̍M������M�� ����T$�B؋J�3������Ė�a�������̍�@�����P���������z����T$������������3��m�������%�����������̋M��H����T$�B��J�3��A����$������������������̋M������T$�B��J�3������P������������������̋M������T$�B��J�3�������|�����������������̋M�鸲���T$�B��J�3���������i���������������̋E�P�����YËT$�B��J�3��~����ԗ�6������������̋E�P�ǚ��YËT$�B�J�3��N���� ��������������̋E�P藚��YËT$�B��J�3������,���������������̋E�P�g���YËT$�B�J�3�������X��������������̋E�P�7���YËT$�B��J�3���������v������������̋E�P����YËT$�B�J�3���������F������������̋E�P�י��YËT$�B��J�3��^����ܘ�������������̋E�P觙��YËT$�B�J�3��.�������������������̋E�P�w���YËT$�B��J�3�������4��������������̋E�P�G���YËT$�B�J�3�������`��������������̋E�P����YËT$�B��J�3���������V������������̋E�P����YËT$�B�J�3��n�������&������������̋M��i���T$�B�J�3��A����������������������̋M���h���M����}����M��� �����T$�B�J�3������� �����������̋E�P�G���YËT$�B��J�3�������L��������������̋E�P����YËT$�B�J�3������x��V������������̋M��x����M����   �L���M����   �L���T$�B��J�3��U����������̋M��8����M����   �zL���M����   �lL���T$�B��J�3������������̋EP�M�Q�CL����ËT$�B��J�3���������������̋M��8����T$�B��J�3�������H��y���������������̋M������T$�B��J�3������t��I���������������̋M�������T$�B��J�3��a����������������������̋M������T$�B��J�3��1����̛�����������������̋M��x����T$�B��J�3������������������������̋M��H����T$�B��J�3�������$�����������������̋M������T$�B��J�3������P��Y���������������̋M�������T$�B��J�3��q����|��)���������������̋M������T$�B��J�3��A�����������������������̋M������T$�B��J�3������Ԝ�����������������̋M��X����T$�B��J�3������� �����������������̋M��(����T$�B��J�3������,��i���������������̋M�������T$�B��J�3������X��9���������������̋M�������T$�B��J�3��Q�������	���������������̋M������T$�B��J�3��!�����������������������̋M��h����T$�B��J�3�������ܝ����������������̋M��d���M���0��F���T$�B�J�3��������n����̋M��hd���M���0��F���M���H��F���M���`�����T$�B�J�3��p����T��(��������������̍M������T$�B܋J�3��A�����������������������̍M��x{���T$�B��J�3�������������������������̋E�P�W���YËT$�B��J�3�������؞�������������̋E�P�'���YËT$�B��J�3��������f������������̋E�P�����YËT$�B��J�3��~����0��6������������̋E�P�ǒ��YËT$�B��J�3��N����\��������������̋E�P藒��YËT$�B��J�3����������������������̋E�P�g���YËT$�B��J�3����������������������̋E�P�7���YËT$�B��J�3���������v������������̋E�P����YËT$�B��J�3��������F������������̋E�P�ב��YËT$�B��J�3��^����8��������������̋M������T$�B��J�3��1����d������������������̋M��x����T$�B��J�3������������������������̋E�P�G���YËT$�B�J�3����������������������̋M������T$�B��J�3��������Y���������������̋M�������T$�B��J�3��q������)���������������̋M������T$�B��J�3��A����@������������������̋E�P臐��YËT$�B��J�3������l���������������̋E�P�W���YËT$�B��J�3����������������������̋M��(����M�������T$�B�J�3������̡�^����̋M�������T$�B��J�3���������9���������������̋E�P�Ǐ��YËT$�B��J�3��N����$��������������̍M��xD���T$��|�����x���3������P������������̋M��&���T$�B�J�3�������|�����������������̋E�P�7���YËT$�B��J�3���������v������������̋E�P����YËT$�B�J�3������Ԣ�F������������̋M��x����T$�B�J�3��a���� �����������������̋M��H����M����}C���M����   ��$���T$�B�J�3������<���������̍M�鸳���T$�B��J�3�������h�����������������̍�p����C���T$������������3���������p������̋E�P����YËT$�B��J�3���������F������������̋EP�׍��YËT$�B��J�3��^������������������̋E�P�M�Q�B����ËT$�B��J�3��(�������������̋E�P�w���YËT$�B�J�3�������D��������������̋M��]���M����=����T$�B�J�3�������x��~����̋M��x]���M��������M���$�����T$�B��J�3���������C���������̋E�P�׌��YËT$�B��J�3��^������������������̋E�P觌��YËT$�B�J�3��.�������������������̋M���\���T$�B��J�3������8�����������������̋M��\���T$�B��J�3�������d�����������������̋E�P����YËT$�B��J�3���������V������������̋E�P����YËT$�B�J�3��n�������&�������������h@jj�E���P�����ËM���,�B���M���<�C���T$�B��J�3����������������������h@jj�E���P�}���ËM���,�/B���M���<��B���T$�B�J�3�������4�������������̋M��xY���T$�B��J�3������`��Y���������������̋E�P����YËT$�B��J�3��n�������&������������̋M��Y���M����E���T$�B�J�3��6������������̍�@����U�����x����j����T$������������3���������������������̋E�P�G���YËT$�B�J�3������� ��������������̋E����   �e���M��>��ËT$�B�J�3������L��H��������������̍M��>���T$��t�����p���3��[����x�����������̋E�P觉��YËT$�B��J�3��.�������������������̋E�P�w���YËT$�B�J�3�������Ч鶿�����������̋M��Ȏ���M����>��h@jj�E��   P�H���ËT$�B��J�3��������f������������̋M��x����M�����=��h@jj�E��   P�����ËT$�B��J�3��^����H��������������̍M��=���T$�B�J�3��1����t�����������������̍M��X=����h����M=����d���P�a���YËT$��L�����H���3���������难���������������̍M��=���M�� =���M���<���M���<���T$��L�����H���3���������K�����������������̍M��<���M��<���M��<���M��<���T$��L�����H���3��C����8��������������������̍M�h<���T$�B��J�3������d��ɽ��������������̋M��8<���M����   �:���T$�B��J�3���������鋽����������������̋M���;���T$�B��J�3������ĩ�Y���������������̋M���c���M����   ��{���T$�B��J�3��c������������������������̋M��c���T$�B��J�3��1����$�����������������̋E�P�w���YËT$�B��J�3�������P�鶼�����������̋E�P�G���YËT$�B�J�3��ο���|�醼�����������̋E�P����YËT$�B��J�3�螿������V������������̋M��h����M����:��h@jj�E��   P������h@jj�E��   P�����ËT$�B��J�3��6����������̍M��h:���M��`:���T$�B؋J�3��	���� ����������̍�x����5:���M��-:���M��%:���M��:���M��:���M��:���E�P�$���YËE�P����YËT$��L�����H���3�蚾���D��R��������̋E�P����YËT$�B�J�3��n�������&������������̍M��l���T$�B��J�3��A����ܫ�����������������̍M��h9���T$�B�J�3��������ɺ��������������̍M�89���T$�B��J�3������4�険��������������̍M��9���T$�B�J�3�豽���`��i���������������̍�P�����8����d�����Y���M���8���T$����������3��e����������̍M��8���T$��L�����H���3��;����Ȭ����������̍�`����e8����P����Z8���T$����������3���������鵹����������̋EP�G���YËT$�B�J�3��μ���(�醹�����������̋E�P����YËT$�B��J�3�螼���T��V������������̍�������7���������7���T$������������3��]������������������̍�P����7����,���������h����o7���T$����������3������ĭ�ʸ���������������̍�8����57���T$����������3��ػ����鐸�����̋M��xD���T$�B�J�3�豻�����i���������������̋M�阜���T$�B��J�3�聻���H��9���������������̋E�P�ǁ��YËT$�B��J�3��N����t��������������̋E�P藁��YËT$�B�J�3���������ַ�����������̋M������M����m����T$�B��J�3������Ԯ鞷���̋M��؛���M����=����M����"/���M���(�7����M���8�\����M���P��5���T$�B�J�3�芺������B��������̋E�P�׀��YËT$�B��J�3��^����T��������������̋M��H����M���魈���M����.���M���(�����M���8������M���P�Q5���M����   �C5���T$�B��J�3������x�餶���������̋E�P�7���YËT$�B�J�3�边���ܯ�v������������̍M��y���T$�B��J�3�葹�����I���������������̍M���x���T$�B��J�3��a����4�����������������̋M���L���T$�B��J�3��1����`�����������������̋M��L���M��� �mx���T$�B�J�3���������鮵���̋M������T$�B��J�3��Ѹ�����鉵��������������̋E�P���YËT$�B��J�3�螸�����V������������̋E�P��~��YËT$�B�J�3��n������&������������̋E�P�~��YËT$�B��J�3��>����D���������������̋E�P�~��YËT$�B�J�3������p��ƴ�����������̋M�������M����-3���M����   ������M����   �1w���M����   �#w���T$�B�J�3�謷������d����������̋M�阘���M�����2���M����   �o����M����   ��v���M����   ��v���T$�B��J�3��L����������������̋M������T$�B��J�3��!����4��ٳ��������������̋M�������M����   �Zv���T$�B�J�3������h�雳����������������̋E�P�'}��YËT$�B��J�3�讶������f������������̋E�P��|��YËT$�B�J�3��~�������6������������̋E�P��|��YËT$�B��J�3��N������������������̋E�P�|��YËT$�B�J�3��������ֲ�����������̋E�P�g|��YËT$�B��J�3������D�馲�����������̋E�P�7|��YËT$�B�J�3�辵���p��v������������̋E�P�|��YËT$�B��J�3�莵������F������������̋E�P��{��YËT$�B�J�3��^����ȳ�������������̋E�P�{��YËT$�B��J�3��.�������������������̋E�P�w{��YËT$�B�J�3������� �鶱�����������̋EP�M�Q�#0����ËT$�B��J�3��ȴ���L�週�����̋E�P�{��YËT$�B��J�3�螴���x��V������������̋M�鈕���T$�B��J�3��q�������)���������������̋E�P�z��YËT$�B�J�3��>����д��������������̋M��(����M����P���M���8�P���M���h�G/���M���x�$���M����   ��#��h@jj�E��   P�Y���ËM����  ������T$�B�J�3�豳������i���������������̋M�阔���M�����O���M���8��O���M���h�.���M���x�|#���M����   �n#��h@jj�E��   P�����ËM����  �8����M����  �Z,���T$�B��J�3������X��˯����������������̋E�P�Wy��YËT$�B��J�3��޲���̵閯�����������̋E�P�'y��YËT$�B�J�3�讲������f������������̋M�阓���M����}���T$�B��J�3��v����,��.����̋M��h����M����M���T$�B��J�3��F����`�������̋E�P�x��YËT$�B��J�3���������֮�����������̋E�P�gx��YËT$�B�J�3��������馮�����������̋M��Ha���M����-���M���8�-���T$�B��J�3�諱������c���������̋M��a���M�����,���M���8��,���T$�B�J�3��k����0��#���������̋M���`���M����,���T$�B��J�3��6����d������̍�H����e,����`����Z,���� ����O,���� ����D,���� ����9,���� ����.,���� ����#,���T$������������3��ư������~����̋E�P�w��YËT$�B��J�3�螰�����V������������̋E�P��v��YËT$�B�J�3��n������&������������̍�0����+����`����+����(���P�v��YËE�P�v��YËT$����������3������\��̬���M��x_���M����=+���T$�B��J�3��������鞬���̋M��H_���M����+���M��� �+���T$�B��J�3�諯���̸�c���������̋M��_���M�����*���T$�B��J�3��v���� ��.����̋E؃��   �e���M�*��ÍM��*���T$�B��J�3��8����4��������̍M�h*���M��`*���T$�B�J�3��	����h����������̋E����   �e���M��(*��ËT$�B܋J�3��Ю�����鈫�������������̍M��)���T$�B�J�3�衮������Y���������������̍M���)���T$�BԋJ�3��q������)���������������̍M��)���T$�B��J�3��A����������������������̍M��h)���T$�B�J�3������D��ɪ��������������̍M��8)���T$�B�J�3������p�陪��������������̋E����   �e���M���(��ËT$�B܋J�3�蠭������X��������������̋E����   �e���M��(��ËT$�B܋J�3��`����Ⱥ���������������̍M��(���M��(���T$�B��J�3��)��������������̍M��X(���M��P(���T$�BЋJ�3�������0�鱩������̍�P����%(���� ����(���������(����0����(���T$������������3�觬���t��_�����̍M���'���T$�B��J�3�聬������9���������������̍M��'���T$�B��J�3��Q����̻�	���������������̋E�P�r��YËT$�B��J�3���������֨�����������̋E�P�gr��YËT$�B�J�3������$�馨�����������̍M�'���T$�B�J�3�������P��y���������������̍M���&����p�����&���M���&���M���&���M���&����d���P��q��YË�d���P��q��YËT$��L�����H���3��L����t������������̍M��x&���T$�B�J�3��!����ؼ�٧��������������̍M������M��@&���T$�B��J�3�������顧������̋M��HZ���T$�B�J�3�������8��y���������������̋E����   �e���M��%��ËT$�B�J�3�耪���d��8��������������̋E�P��p��YËT$�B�J�3��N�������������������̋E�P�p��YËT$�B��J�3���������֦�����������̋M��xY���M����i���M����   �/%���T$�B��J�3��ة�����鐦�����̋M��8Y���M����]i���T$�B�J�3�覩���,��^����̋M��Y���M����-i���T$�B�J�3��v����`��.����̋M���X���M�����h���T$�B��J�3��F������������̍������u$���������j$���T$������������3������Ⱦ�ť����������̍M��8$���E����   �e���M�� $��ËT$��L�����H���3��¨������z����������������̍M���#����p�����#���M���#���M���#���M���#���M��#���M��#���T$��L�����H���3��X���� ��������̍�l�����t���T$��d�����`���3��(�������������̋E�P�wn��YËT$�B��J�3���������鶤�����������̋E�P�Gn��YËT$�B�J�3��Χ���ܿ醤�����������̍�������"����(����Jg����������"���T$������������3�肧�����:����������������̍������"����(�����f���������"���T$������������3��2����T������������������̍M��X"���M��P"���E�P�gm��YËE�P�\m��YÍM��2"���M��*"���M��""���M��"���T$��L�����H���3�车���x��u�����������̍�������!���T$������������3�舦������@������̍M���B����P����!���T$����������3��P��������������������̍� ����u!����<����B���������_!���������������@����I!���T$������������3������<�餢���������̍�<����uT���T$��4�����0���3�踥������p������̍M��� ���M��� ���T$�B��J�3�艥������A�������̍M�� ���M�� ���T$�B��J�3��Y��������������̋E�P�k��YËT$�B��J�3��.����$��������������̍M��Hd���T$�B�J�3������P�鹡��������������̋E����   �e���M� ��ËT$�B�J�3�������|��x��������������̍M��s���M������T$�B��J�3�艤������A�������̋M��8;���T$�B��J�3��a����������������������̋M��;���M����c���T$�B��J�3��&������ޠ���̋E�P�wj��YËT$�B��J�3�������<�鶠�����������̋E�P�Gj��YËT$�B�J�3��Σ���h�醠�����������̋M��x:���M����c���M����   ��b���M����   ��b���M����   ��b���T$�B��J�3��l�������$����������̋M��:���M����b���M����   �b���M����   �b���M����   �b���M����   �ub���T$�B��J�3���������鶟�����������̋M�� ���M����   銿���T$�B܋J�3��â���<��{�����������������̋M��H ���T$�B��J�3�葢���h��I���������������̋E�P��h��YËT$�B��J�3��^�������������������̋E�P�h��YËT$�B�J�3��.�������������������̋E�P�wh��YËT$�B��J�3���������鶞�����������̋E�P�Gh��YËT$�B�J�3��Ρ����醞�����������̋M��x8���M����a���T$�B��J�3�薡���L��N����̋M��H8���M�����`���T$�B��J�3��f�����������̋M��8����T$�B��J�3��A�����������������������̋E�P�g��YËT$�B�J�3���������Ɲ�����������̋E�P�Wg��YËT$�B�J�3��ޠ����閝�����������̋E�P�'g��YËT$�B�J�3�讠���0��f������������̍M��_���T$�B�J�3�聠���\��9���������������̋M��H����T$�B��J�3��Q�������	���������������̋E�P�f��YËT$�B��J�3���������֜�����������̋E�P�gf��YËT$�B��J�3��������馜�����������̋E�P�7f��YËT$�B��J�3�辟�����v������������̋M����e����T$�B��J�3�莟���8��F������������̍�(����_���T$����������3��X����d��������̍M�����T$����������3��+����������������̍�X����;����@���������T$��8�����4���3��������饛����������̍M�����T$�B��J�3����������y���������������̍M������T$��L�����H���3�苞�����C���������̍M���l���T$�BȋJ�3��a����H�����������������̍M�����M�����T$�B��J�3��)����|���������̋M��j���T$�B��J�3��������鹚��������������̋M��hj���T$�B��J�3��ѝ�����鉚��������������̍M�����T$�B��J�3�衝��� ��Y���������������̍M�����T$�B�J�3��q����,��)���������������̍M�����T$�B�J�3��A����X������������������̍�X����9����T������   ��T�����M�G��ËT$��T�����P���3��������顙������̍M����T$�B��J�3����������y���������������̍�\���������l����i���T$��\�����X���3��}�������5�����������̍�8�����h����(�������T$����������3��=���� ��������������̍M�h���M��h���M����   �R���T$�B��J�3�������\�鳘��������̍M��(���T$�B�J�3��ћ�����鉘��������������̋M��8h���M����   �����T$�B��J�3�蓛������K�����������������̍�p�������T$����������3��X�������������̍�d�������������z���������o���T$��h�����d���3������$��ʗ���������������̋M��8���T$�B��J�3������P�陗��������������̋�x������   ��x�����M����ËT$��t�����p���3�蔚���|��L����M������M������T$������������3��c������������������������̋M���H�u����M����   �����T$�B��J�3�� �������ؖ�������������̋E�P�g`��YËE�P�\`��YËT$�BԋJ�3�������雖����������������̋M�������T$�B��J�3�讙���D��f������������̋M��������T$�B��J�3��~����p��6������������̍���������T$��L�����H���3��H������� ������̋M�������T$�B�J�3��!�������ٕ��������������̋E�P�g_��YËT$�B��J�3��������馕�����������̋E�P�7_��YËT$�B�J�3�辘��� ��v������������̍M������T$�BԋJ�3�葘���L��I���������������̍�(��������8��������H�������T$������������3��B������������������������̋�����P�^��YËT$������������3��������齔��̍M��8���M��0���T$�BԋJ�3��ٗ�����鑔������̍M�����M�� ���T$�BЋJ�3�詗�����a�������̍M�������h��������T$��L�����H���3��p������J�3��c����P�������������������̍M������x����}���T$��p�����l���3�� ������J�3���������˓����������������̍M��8���E�P�O]��YËE�P�D]��YËE�P�9]��YÍ�d���������x��������T$��@�����<���3�褖������\����M������M������M������M������T$�B��J�3��i������!�������̋EP�M�Q�����ËT$�B��J�3��8����H��������̍M��h���T$�B��J�3������t��ɒ��������������̋E�P�W\��YËT$�B��J�3��ޕ�����閒�����������̋E�P�'\��YËT$�B��J�3�讕������f������������̋M��X,���M����ͬ���T$�B�J�3��v���� ��.����̋M��(,���M���靬���T$�B��J�3��F����4�������̋EP�M�Q�s����ËT$�B��J�3������`��Б�����̋E�P�g[��YËT$�B��J�3��������馑�����������̋E�P�7[��YËT$�B�J�3�辔������v������������̋E�P�M�Q������ËT$�B�J�3�舔������@������̋M��8����T$�B��J�3��a���������������������̋M�������M����   �z����T$�B�J�3��#����D��ې����������������̋M������T$�B��J�3������p�驐��������������̋E�P�7Z��YËT$�B��J�3�输������v������������̋E�P�Z��YËT$�B�J�3�莓������F������������̍������Ŷ���T$������������3��X�������������̋M��� �R���M���$�R���M���(�R���M���,�R���M���0�yR���M���4�nR���M���8�cR���M���<�XR���M���@�MR���M���D�BR���M���H�7R���T$�B��J�3���������x��������������̋M��h)���M�����Q���T$�B�J�3�膒������>����̋E�P��X��YËT$�B��J�3��^�������������������̋M��)���M����Q���M����Q���M���@�#���T$�B�J�3��������Ȏ�������������̋E�P�WX��YËT$�B�J�3��ޑ���@�閎���M������T$�B�J�3�軑���l��s����M�鿴���T$�B�J�3�蘑������P����T$�B�J�3��}����@��5������������j j j ��8�=������������������h�   h�   h�   ��8�g=���������j j j ��8�P=������������������h�   h�   h�   ��8�'=���������h��[���Y�����V�   ����`9^��������������V�   �����h9^��������������V�   �������p9^������������V�   �e���x9^��������������V�   �E���|9^��������������V�   �%������9^�����������̡P9h43h03h$3�������]#�����   �h �^���Y��������h0�K���Y�����h�8h0�h�h$3h�8��9��*��hp����Y��h�8hph��h�8h�8��:�*��h�����Y��h(9h �h0�h�8h9��;�*��h�踣��Y��h�;h �h@�h$3h�;��<�]*��h�舣��Y��h��{���Y�����hTCh 'h�%hHCh8C�H>�*��h��H���Y��hEj j hEhHC�8?��)��h�����Y��������hUh�"hPhEh U�8@�)��h�����Y��V� A腰��h��Т����^�������V��A�Ű��h 谢����^�������hDUh��h`�hEh0U��A�M)��h�x���Y��h|Uh �h �hEhlU��B�)��h �H���Y��h�Uh��h��hEh�U��C��(��h0����Y��h�Uh`�h��h�8h�U��D�(��h@����Y��h8Vh��h��h�8hV��E�(��hP踡��Y��h�^hP5hPHhEh�^��F�](��h`舡��Y��h_h�6h 6hEh_�pG�-(��hp�X���Y��hd_hpOhLh�8hD_�XH��'��h��(���Y��h�_h09h@8h�8h�_�@I��'��h������Y��hih�h �hih�h�0J�'��h��Ƞ��Y��hTih��h��h�8h@i�K�m'��h�蘠��Y��hh�h�	h��h\�hL��L�='��h��h���Y��h��h
h �h��h��� M�'��h��8���Y��h�hPh0�h��hԪ��M��&��h�����Y��h�h�h��hEh���N�&��h��؟��Y��hX�h�h��hH�h<���O�}&��h 訟��Y��h��h hhEh����P�M&��h�x���Y��hP�h� h�hEh\���Q�&��h �H���Y��h|�hP�h0�hEhp���R��%��h0����Y������U����hS���������������h��h09h�=h$3hx���S�%��h@�Ȟ��Y��h��h`"h`0h$3h���hT�m%��hP蘞��Y��h��h &hP1h$3h���PU�=%��h`�h���Y��h,�huh thEh ��@V�%��hp�8���Y��� 5���\$�(W�@'�\$�X��$�����������j��;��Pj�@W�L=���HW���PW�I����'�XWh��P<�pW    �`W�tW   �p&�hW蜝��Y������hD&h�1	h�0	h�8h$&��W�=$��h��h���Y��h@,h0�
h��
hHCh,,��X�$��h��8���Y��U�������tSVW���T$�L$P���\$�$���������T$�L$h�\$�����$�ܼ������T$�T$��$�   �$��込���hY��������Y������Y�޻����Y�Ի����Y�z���VWS�hY譓��h�舜����_^[��]����������U�������tSVW���\$�L$P���T$�$�9�������T$��L$h���\$�$��������T$��$�   �T$���$�������Y���2���� Z�(����Z�����0Z�����HZ����VWS��Y����h��ț����_^[��]����������U�������tSVW���T$�L$P�\$���$�y�������\$��L$h���T$�$�\�������T$�T$��$�   �$���>����hZ���r�����Z�h�����Z�^�����Z�T�����Z�����VWS�hZ�-���h�������_^[��]����������VW�    �hY��Zh���ؚ����_^��������������hd2h@�
h��
hihT2��c�m!��h�蘚��Y��hx4hph�hihh4�pd�=!��h �h���Y��h�8h�Qh�Phih�8�`e�!��h�8���Y��h�<h��hP�hHChp<�Pf�� ��h ����Y��h\@j j h$3h�8�Hg� ��h0�ޙ��Y��������h�@h@�h �h�8h�@�0h�} ��h@訙��Y��h�@h��h��h�8h�@�i�M ��hP�x���Y��hAh �h@�h$3h�@� j� ��h`�H���Y������T$��j�\$���$��������T$�\$� k�0'�$�����hp�����Y���������hOhP:h@gh�8h O�Hk���h��Ș��Y��hLOh�;h0hh�8h8O�0l�m��h�蘘��Y��h�Oj j hEhtO�m�C��h��n���Y��������h�Oh ih��htOh�O� n���h��8���Y��h�Oh�=h��htOh�O��n����h�����Y��h<Ph >h��htOh$P��o���h��ؗ��Y��htPh�>h��htOhdP��p�}��h�託��Y��h�Ph�>h��htOh�P��q�M��h��x���Y��h�Ph@h ?hEh�P��r���h �H���Y��hQh�@h��htOhQ�ps����h����Y��h`Qh Xh Wh�8hDQ�Xt���h ����Y��h�Qhpehpdh�8h�Q�@u���h0踖��Y��h�Sh��h��h$3h�S�0v�]��h@舖��Y��h Zh0�h��h$3hZ� w�-��hP�X���Y��h�^h@�h@�h�8h�^�x����h`�(���Y��h _hp�hp�h$3h�^� y����hp�����Y��h4_h �h�hEh(_��y���h��ȕ��Y��h�_h�h`h$3h�_��z�m��h�蘕��Y��hah�h@hH�h�`��{�=��h��h���Y��h,bhp+hP*hihH���|���h��8���Y��h�dhPNh0Mhih�d��}����h�����Y��h8ehOh�Nh�dh e��~���h��ؔ��Y��h\fj j hEhi�����h�讔��Y��������h8gh��hЊhEh(g�p��M��h��x���Y������T$�X��T$�$�F���������hhhp�h��hEhh�x�����h �(���Y��h�lj j hEh�l�������h�����Y��������h mh��h��h�lhm�p����h �ȓ��Y��h\mh��hЭh�lhHm�X��m��h0蘓��Y��h�mh0�h�h�lh�m�@��=��h@�h���Y��h�mh��h��h�lh�m�(����hP�8���Y��hnh�h �h�lh�m������h`����Y��hDnh�h�h\�h,n������hp�ؒ��Y��h�nhP�h`�hEhln����}��h�訒��Y��h sh �h@�hEh�r�Љ�M��h��x���Y��h8sh��h`�hEh(s������h��H���Y��h�sh��h �hEh�s�������h�����Y��h�uh �h0�hHCh�u������h�����Y��h�wh h hHCh��������h�踑��Y��hzh�1hp0hHCh�y�x��]��h�舑��Y��h�}h0LhKhHChx}�h��-��h��X���Y��h�}j h lhx}h�}�P�� ��h �+���Y�����hX~j j h$3hE�@�����h�����Y��������h�h�vhp{h$3h��0����h �Ȑ��Y��h��h��h�h�8h܀� ��m��h0蘐��Y��h$�h��hЊh$3h����=��h@�h���Y��h�j j h$3h�� ����hP�>���Y��������hL�h@�h��h�h8�������h`����Y��h��h �h�h�ht��Ж���hp�؏��Y��hĄh �hP�h8�h������}��h�訏��Y��h�h �h��h�8h������M��h��x���Y��h��h`�h`�h�8hl�������h��H���Y��hĜh`�h��h$3h���������h�����Y��h��h��h��h$3h��p����h�����Y��h|�h�%h�!h$3hl��`����h�踎��Y�̃=�8 uK��8��t��8�Q<P�B�Ѓ���8    ��8��tV������V�Z@������8    ^����������������������������3���9��9��9��9��9��9��9��9��9��9��9������̹�9����������̹�:���������̹�;���������̹�<�������������������������̹H>�v��������̹8?�f��������̹8@�V����������������������������������������̹�A�&��������̹�B���������̹�C���������̹�D����������̹�E����������̹�F����������̹pG����������̹XH���������̹@I���������̹0J���������̹K���������̹L�v��������̹ M�f��������̹�M�V��������̹�N�F��������̹�O�6��������̹�P�&��������̹�Q���������̹�R���������̹�S����������̹hT����������̹PU����������̹@V����������̹PW��6�������̹�W���������̹�X�������������������������������������������������������������������������̹�c�F��������̹pd�6��������̹`e�&��������̹Pf���������̹Hg���������̹0h����������̹i����������̹ j��������������������������̹Hk���������̹0l���������̹m���������̹ n���������̹�n�v��������̹�o�f��������̹�p�V��������̹�q�F��������̹�r�6��������̹ps�&��������̹Xt���������̹@u���������̹0v����������̹ w����������̹x����������̹ y����������̹�y���������̹�z���������̹�{���������̹�|���������̹�}�v��������̹�~�f��������̹��V��������̹p��F��������̹x��6��������̹���&��������̹p����������̹X����������̹@�����������̹(�����������̹�����������̹������������̹�����������̹Љ���������̹�����������̹�����������̹���v��������̹���f��������̹x��V��������̹h��F��������̹P��6��������̹@��&��������̹0����������̹ ����������̹�����������̹ �����������̹�����������̹Ж����������̹�����������̹�����������̹�����������̹�����������̹p��v��������̹`��f���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ��     ��     Z� f� z� �� �� �� �� �� � � "� 2� >� P� `� n� �� �� �� �� �� �� �� �� � � $� 0� H� `� j� v� �� �� �� �� �� �� �� �� D� 
� $� <� V� l� �� �� �� �� �� �� �� �  � 0� F� V� d� v� �� �� �� �� �� �� �� � � ,� B� R� .� � � �� �� �� �� ��     ��     p� |�         ��������� �@�`��������� �0�`������� �0�`������� �0�`������� �P������� @ p � �  0`���@p�@ ����@p�� 0���@p�� 	0	`	�	�	�	 
P
�
�
�
@p��  P���@p�� 0`��� P���@p�� 0`�        
������.�        �U�                �YU       k    �  � bad allocation  ���� � LP  L�K�K�K%   +   c:\program files\maxon\cinema 4d r12\plugins\rhinoio\source\register.cpp    ?name=  &organization=  &street=    &city=  &country=   &c4dserial= ���ư>H�0 ֌         �f@-DT�!	@              �?�������������      �?   �MbP?3D Geometry File Format  ��� �� �  � H� � Ф 0� @� ��P� ��  �  � ع�� Ф 0� @�  �� Ф 0� @�     c:\program files\maxon\cinema 4d r12\resource\_api\ge_dynamicarray.h    ���� * @r`rpr�9 Pr�r�r�r�r�rs�+  s�r�r�,  b rhino_docs_us.html  file:// #import help    rhino_docs_ .html   c:\program files\maxon\cinema 4d r12\plugins\rhinoio\source\rhinoloader.cpp        @R��?{�G�z�?     @�@ - Red   - Green     - Blue     es-8R��?:�0�yE>Frhinoimport    ��P@� D�P@� vector<T> too long  
        @P�Rhino Import Error: Selection Include List not found!         �      �?      �?      @      B@ ���\�B  ��~5�B   \]աAo��ʡ�?UUUUUU�?�q�q�?����MbP?���ư>    ��.A     @�@      Y@      $@�������?rb      ���ư>c:\program files\maxon\cinema 4d r12\plugins\rhinoio\source\rhino.h     л�� �� @r`rpr`� Pr�r�r�r�r�rs s s�r�rP� #export     c:\program files\maxon\cinema 4d r12\plugins\rhinoio\source\rhinosaver.cpp  Frhinoexport    3dm       >@      N@$�P@� map/set<T> too long invalid map/set<T> iterator Rhino Export: Major point sort error!       Rhino Export: Mesh self test failed, not inserted into the document!    Rhino Export: Writing the model to file unsuccessful!   -> other spline (   )   Rhino Export: Polyline invalid! autschn!              2@t��*�*��rhinoi  %08X    c:\program files\maxon\cinema 4d r12\plugins\rhinoio\source\serial.cpp  ���8c:\program files\maxon\cinema 4d r12\resource\_api\c4d_resource.cpp #   M_EDITOR    <��Kres c:\program files\maxon\cinema 4d r12\resource\_api\c4d_general.h    %s         -DT�!��-DT�!�?-DT�!@�h㈵��>       @      �A      �A
ףp=
�?       �
ףp=
�?      @c:\program files\maxon\cinema 4d r12\resource\_api\c4d_file.cpp ����̽�    c:\program files\maxon\cinema 4d r12\resource\_api\c4d_baseobject.cpp   �P�`SpS�S�S�S�S�S�'`�P�`SpS�S�S�S�S�S�T����0d@d�d�dPd�d�d�d e�ec:\program files\maxon\cinema 4d r12\resource\_api\c4d_gui.cpp  ��P�`SpS�S�S�S�S�S�h@�P�`SpS�S�S�S�S�S�pq q0q@qPq`qpq`��q�q�q�qProgress Thread 0%  ~   ����Б��c:\program files\maxon\cinema 4d r12\resource\_api\c4d_basebitmap.cpp   c:\program files\maxon\cinema 4d r12\resource\_api\c4d_pmain.cpp        c:\program files\maxon\cinema 4d r12\resource\_api\c4d_libs\lib_ngon.cpp        c:\program files\maxon\cinema 4d r12\resource\_api\c4d_basetime.cpp      �Ngm��C   ����A  4&�k�  4&�kC�����W������    c:\program files\maxon\cinema 4d r12\resource\_api\c4d_gv\ge_mtools.cpp 4� |����`                �������������������YLN��i�Gl�<�����H�����O~F:��K�M�KVR���_Q`��A���/��@#/��NI��o�|�C�j�G��|Wy��cS)?�D��D��~'9����EN�g��پR����W�%F�����0�.\opennurbs_object.cpp  ON__dblinithelper   CPU has unexpected bit pattern in double 2.0.   ON__fltinithelper   CPU has unexpected bit pattern in float 2.0f.      @���W�' ���`����W� �ON_Object::ClassId() FAILED
    class uuid:     class name: %s
 unknown ON_ClassId::ON_ClassId() - class uuid is nill.  ON_ClassId::ON_ClassId() - class uuid already in use.   ON_ClassId::ON_ClassId() - missing baseclass name.  ON_ClassId::ON_ClassId() - class name already in use.   ON_ClassId::ON_ClassId() - class name already in use.  Will append number to make it unique.    ON_ClassId::ConstructorHelper   ON_ClassId::ON_ClassId() - missing class name   ON_Object::AttachUserData       ON_Object::AttachUserData() - attempt to attach invalid UnknownUserData.    ON_Object   0   60B5DBBD-E660-11d3-BFE4-0010830122F0    CRC List: %08x, %08x, %08x, %08x, %08x, %08x, %08x, %08x
   Last Modified Time: %u (seconds since January 1, 1970, UCT)
    Size: %llu bytes
   zero (not set)
 Checksum:   .\opennurbs_string.cpp  ON_String::Empty    ON_String::Empty() encountered invalid header - fixed.      p?     �o@      �<L    ;.\opennurbs_xform.cpp   ON_Xform::Rotation  sin_angle and cos_angle are both zero.      �������?�    P>   ����?      ��3�����-C��6?                            	   
                                              	   
                  0123456789abcdef                                                            Layer name is empty.
   L a y e r   E x t e n s i o n s     X���W q �r�`����W� �    ���q��p� �r��r�r�s�t�W� ��u�u�S a v e d   L a y e r   S e t t i n g s     ,� ��	����default material index = %d
    plot color rgb =    display color rgb =     picking = %s
   unlocked    locked  display = %s
   hidden  visible name = "%ls"
   index = %d
     .\opennurbs_layer.cpp   ON_Layer::Read  ON_Layer::Read() encountered a layer written by future code.        t��p��P� �r��� �p��W� ��p����� � �@����Pk��� 0l x`��x {`l� �ON_Layer    95809813-E985-11d3-BFE5-0010830122F0    ON__LayerExtensions ON_UserData 3E4904E6-E930-4fbc-AA42-EBD407AEFE3B    ON__LayerSettingsUserData   BFB63C09-4BC7-4727-89BB-7CC754118200    �7��1!�O��U$�������J��A��~�.\opennurbs_3dm_attributes.cpp  ON_3dmObjectAttributes::ReadV5Helper    Bug in ON_3dmObjectAttributes::ReadV5Helper or WriteV5Helper    Object rendering attributes are not valid.
 Object id is nil - this is not valid.
  X�`��#	@��0���P���@/%d  ,%d groups:     material source = %s
   layer material  object material parent material object material index = %d
 object layer index = %d
    object mode = %s
   normal  object uuid =   object name = "%ls"
    ���p0 ��00�0��� � P���0�� ���W� �ON_3dmObjectAttributes  A828C015-09F5-477c-8665-F0482F5D6996                 �      �=%.17g to %.17g, %.17g to %.17g, %.17g to %.17g
 not valid   Bounding box:       ��&�.>�-���q=9�R�Fߑ?      P=      �>      �  CV      NULL cv array
    Control Points  %d %s points
  index               value
   non-rational    rational    Knot Vector ( %d knots )
   ON_NurbsCurve dim = %d is_rat = %d
        order = %d cv_count = %d
    cv[%d*cv_stride + %d] = %g is not valid.
       cv_stride = %d and cv_size = %d (cv_stride must be >= cv_size).
    cv_size = %d (must be >= 1).
   cv_count = %d (must be >= 2).
  cv pointer is null.
    ON_NurbsCurve is a line with no length.
    ON_NurbsCurve.m_cv has zero weights for CV[%d].
    ON_NurbsCurve.m_cv has zero weights for CV[%d],...,CV[%d].
 ON_NurbsCurve.m_cv has a zero denominator in the parameter interval [%g,%g].
   ON_NurbsCurve.m_cv[] is not valid.
 ON_NurbsCurve.m_knot[] is not a valid knot vector.
 ON_NurbsCurve.m_knot is NULL.
  ON_NurbsCurve.m_cv is NULL.
    ON_NurbsCurve.m_cv_stride = %d (should be >= %d).
  ON_NurbsCurve.m_cv_count = %d (should be >= m_order=%d).
   ON_NurbsCurve.m_order = %d (should be >= 2).
   ON_NurbsCurve.m_dim = %d (should be > 0).
      �c
   9      0@.\opennurbs_nurbscurve.cpp      |���P&�3 ������0�p���p�� �p10�P]@@�0/0/ ��W��p0p��0����3������= ��  �5��>�� �0�n`y������ P p%�� ^
 ^
    )\���(�?{�G�z���������?ffffff�?�������?ON_NurbsCurve::ON_InsertKnot(): knot_multiplicity < 1 or knot_multiplicity > degree.    ON_InsertKnot(): knot_value not in NURBS curve domain.  ON_InsertKnot(): knot_value = t1 and 1 < knot_multiplicity < degree.    ON_NurbsCurve::InsertKnot       ON_InsertKnot(): knot_value = t0 and 1 < knot_multiplicity < degree.    ON_NurbsCurve::Trim ON_NurbsCurve::Trim() - right end de Boor algorithm failed. ON_NurbsCurve   ON_Curve    4ED7D4DD-E947-11d3-BFE5-0010830122F0        D� ;�W I ����;���p�� �����P]@�p�
�
�n�W��p0p�����]
 !	�<����=���= ` !	@c�>0x��P?�W`IPh���A�A���@G�]
�]
�WHH    UUUUUU�?UUUUUU�?     �?empty span. .\opennurbs_curve.cpp   ON_NurbsCurve::SpanIsLinear span_index out of range.        �������?X� ]��<���`~��<�ON_Geometry 4ED7D4D7-E947-11d3-BFE5-0010830122F0    ¦���a�E���~��       ����?     �?  ��false   true        �D�JW�?�������?.\opennurbs_mesh.cpp    ON_MeshParameters::Write    ON_MeshParameters::Read() - m_face_type out of bounds.      �D�JW�?ON_MeshParameters::Read �u �<�7~Y���n���p�� � @�� ����0�� � ��� r@��
�
�n�W��q<����� � @� �p����@�� � ��� r@��
�
�n�W���q��� ��� ��P�p������� � �@� r@��
�
�n�W���qm_mesh=%08x, m_mesh_fi=%d
  mesh xform:
    mapping crc: %08x
  mapping id:     Texture/color coordinates tag:
 O N _ M e s h   d o u b l e   p r e c i s i o n   v e r t i c e s       ����`� � �r�������@��W� �@����C u s t o m   R e n d e r   M e s h   P a r a m e t e r s   ,��		`V`���t���@�����0���<����0��:0�L�г0��:0��� ����8�7��p�� 	 ���$������0�l�P�� �@����0��:0���p	0��:0�D�@� ����(ON_Mesh::Read - compressed vertex color buffer size is wrong.   ON_Mesh::Read - compressed vertex curvature buffer size is wrong.       ON_Mesh::Read - compressed texture coordinate buffer size is wrong. ON_Mesh::Read - compressed vertex normal buffer size is wrong.  ON_Mesh::Read_2 ON_Mesh::Read - compressed vertex point buffer size is wrong.   ����`V`����������?    _�B@��x�D)
  ,   (   m_top_vi = %d (should have 0 <= m_top_vi < %d)
     m_mesh_vi=%d is not in m_top->m_topv[m_top_vi=%d].m_vi[] array.
    m_top_vi = %d and MeshTopology()=NULL
  m_mesh_vi = -1 and m_top_vi = -1
   m_mesh_vi = %d (should have 0 <= m_mesh_vi < %d)
   m_mesh = NULL
  m_top_ei = %d (should have 0 <= m_top_ei < %d)
 m_mesh_fi = %d (should have 0 <= m_mesh_fi < %d)
   ���� �p� �r�@�`� ����W� �������Location:   m_mesh=%08x m_mesh_vi=%d m_top_vi=%d
   m_fCRC != ON_MeshDoubleVertices::FloatCRC(mesh->m_V)    m_fcount != mesh->m_V.Count()   0 = ON_Mesh::Cast( Owner() )    m_dCRC != DoubleCRC()   m_dcount != m_dV.Count()    ON_MeshDoubleVertices::Archive  m_fcount != m_dcount     to     m_mesh=%08x, m_top_ei=%d
   ON_Mesh.m_F[%d] has degenerate double precision vertex locations.
  ON_Mesh.m_F[%d].vi[] has invalid vertex indices.
   Double precision vertices appear to be ok but are not marked as valid
  Single and double precision vertices are not synchronized.
 ON_Mesh.m_vbox is not finite.  Check for invalid vertices
  ON_Mesh.m_N[%d] is not a unit vector (length = %g).
    Single precision vertices appear to be ok but are not marked as valid
  =
ףp=�?��Q���?ON_Mesh.m_S.Count() = %d (should be 0 or %d=vertex_count).
 ON_Mesh.m_T.Count() = %d (should be 0 or %d=vertex_count).
 ON_Mesh.m_N.Count() = %d (should be 0 or %d=vertex_count).
 ON_Mesh.m_V.Count() < 3 (should be at least 3).
    ON_Mesh.m_F.Count() < 1 (should be at least 1).
    m_FN[%d] = (%g,%g,%g)
  %d mesh face normals:
  m_F[%d].vi = (%d,%d,%d,%d)
 m_F[%d].vi = (%d,%d,%d)
    %d mesh faces:
 m_S[%d] = (%g,%g)
  %d mesh vertex surface parameters:
 m_T[%d] = (%g,%g)
  %d mesh vertex texture coordinates:
    m_N[%d] = (%g,%g,%g)
   %d mesh vertex normals:
    m_V[%d] = (%g,%g,%g)
   m_V[%d] = (%.17g,%.17g,%.17g) D = (%.17g,%.17g,%.17g)
  ...
    %d mesh vertices:
  m_Ttag:
    m_srf_scale: %g,%g
 m_srf_domain: (%g,%g)x(%g,%g)
  m_packed_tex_domain: (%g,%g)x(%g,%g)
   m_packed_tex_rotate: %s
    m_Ctag:
    vertex colors:    %s
   vertex kappa:     %s
   tex coords:       %s
   srf parameters:   %s
   face normals:     %s
   vertex normals:   %s
   double precision: %s
   ON_Mesh: vertex count = %d  facet count = %d
          @ON_Mesh::Transform      ON_Mesh::Transform() cannot apply this transform to curvatures.
        $� @"#p� �@�`��� �� ��0� ���P�@P0/0/��W��p`�ON_Mesh::Read   ON_Mesh::Read - surface parameter buffer size is wrong. ON_Mesh 4ED7D4E4-E947-11d3-BFE5-0010830122F0    ON_MeshVertexRef    C547B4BD-BDCD-49b6-A983-0C4A7F02E31A    ON_MeshEdgeRef  ED727872-463A-4424-851F-9EC02CB0F155    ON_MeshFaceRef  4F529AA5-EF8D-4c25-BCBB-162D510AA280    ON_MeshDoubleVertices   17F24E75-21BE-4a7b-9F3D-7F85225247E3    ON_PerObjectMeshParameters  B5628CA9-82C4-4CAE-9883-487B3E4AB28B    ���ư>ON_InstanceDefinition.m_idef_update_type value is invalid.
     ON_InstanceDefinition is linked_and_embedded_def but m_idef_layer_style is not zero.
   ON_InstanceDefinition is linked_def but m_idef_layer_style is not 1 or 2.
      ON_InstanceDefinition is linked or embedded but m_source_archive_checksum is zero.
     ON_InstanceDefinition is linked or embedded but m_source_archive is empty.
     ON_InstanceDefinition.m_idef_update_type = obsolete "embedded_idef". Use "static_def" or "linked_and_embedded_def".
    ON_InstanceDefinition is static but m_idef_layer_style is not zero.
    ON_InstanceDefinition is static but m_source_archive_checksum is set.
  ON_InstanceDefinition is static but m_source_archive is not empty.
 ON_InstanceDefinition has invalid bounding box.
    ON_InstanceDefinition has nil uuid.
    .\opennurbs_instance.cpp    ON_InstanceDefinition::IdefUpdateType       Using obsolete ON_InstanceDefinition::embedded_def value - fix code.    t�*p6@7 �+�`�0,�, -� � �- r@�.0/0/�n�W��pqON_InstanceRef has singular m_xform.
   ON_InstanceRef has nil m_instance_definition_uuid.
     L i n k e d   I n s t a n c e   D e f i n i t i o n   L a y e r   S e t t i n g s       ���/�80: 01�P1p1�12�W� ��2�2�    L i n k e d   I n s t a n c e   D e f i n i t i o n   A l t e r n a t e   P a t h   �@<0��:0�\�=��<�    ��0&�H@I @&�?�5��B`I�(@ � � ) r@��
�
�n�W��pqContains: %d objects
   none.
  Archive     Update depth: %d
   Alternate archive: "%ls" (%s)
  "%ls" (%s)
 absolute    relative    Source archive:     URL tag: "%ls"
 URL: "%ls"
 Description: "%ls"
 Id:     not valid   linked - definition from source archive.    embedded and linked - definition from source archive.   OBSOLETE embedded_def with empty source archive - should be static_def. OBSOLETE embedded_def with non-empty source archive - should be linked_and_embedded_def.    embedded.   Type:   Name: "%ls"
    ��@/�N�L �r�P/`7�7`G�W� �`/08�ON_InstanceDefinition   26F8BFF6-2618-417f-A158-153D64A94989    ON_InstanceRef  F9CFB638-B9D4-4340-87E3-C56E7865D96A    ON__IDefLayerSettingsUserData   11EE2C1F-F90D-4C6A-A7CD-EC8532E1E32D    ON__IDefAlternativePathUserData F42D9671-21EB-4692-9B9A-BC3507FF28F5              �?      �=polycurve.Segment(%d).Domain() does not match polycurve.SegmentDomain(%d).
 polycurve.SegmentCurve(%d) is not closed.
  polycurve.SegmentCurve(%d) is null.
    polycurve.BoundingBox() z values are not both 0.0.
 polycurve.BoundingBox() is not valid.
  polycurve dimension = %d (should be 2).
    polycurve has < 1 segments.
    D��^��н �`�pd�dpe�f�h��` � n0p@s�
�
�n��0��p�B����@�0�P��� ������`�p��� ��@� ���@�`�Ф�����Я � ���%s
 m_path has zero length. m_path has zero length <= ON_Extrusion::m_path_length_min.  m_path has zero direction.  m_t does not satisfy 0<=m_t[0]<m_t[1]<=1    m_N[1].z is too small (<=ON_Extrusion::m_Nz_min) or negative    m_N[1] is not a unit vector.    m_N[0].z is too small (<=ON_Extrusion::m_Nz_min) or negative    m_N[0] is not a unit vector.    m_up is not perpendicular to m_path.    m_up is not a unit vector.  m_profile is not valid.     m_profile_count > 1 but a m_profile_count->SegmentCurve() is not closed.        m_profile_count > 1 but a m_profile_count->SegmentCurve() is null.  m_path is not valid.    m_profile is not a valid ON_PolyCurve.      m_profile_count > 1 but m_profile_count != m_profile->SegmentCount().   m_profile_count > 1 but m_profile is not an ON_PolyCurve.   m_profile is NULL.  m_profile_count < 1.    u    �>      �?m_mesh[%d] = 
  m_mesh[%d] = null
  no cached meshes
   ON_DisplayMeshCache user data
  Cached meshes   .\opennurbs_beam.cpp         @�>��� �� @��������P��W� �к�0�%s %s mesh: %d polygons
    Quality Fast    Custom  preview mesh    analysis mesh   render mesh NULL    Profile:
   Profile Count: %d
  m_bTransposed = %d
 m_path_domain = (%.17g, %.17g)
 ,   m_N[] = (   m_bHaveN[] = (%d, %d)
  m_bCap[] = (%d, %d)
    Up:         Path:   ON_Extrusion: 
 $�����0�p�extrusion has no profile curve. corrupt extrusion cannot produce a brep form.   Failed to add caps to extrusion brep form.  Corrupt extrusion cannot produce brep form. Corrupt profile domain. unable to duplicate profile segment.    null profile segment.   Unable to get allocate brep.    Unable to get top cap location. Unable to get bottom cap location.  ON_Extrusion::BrepForm  extrusion direction is zero.    ON_Extrusion    ON_Surface  36F53175-72B8-4d47-BF1F-B4E6FC24F4B9    ON_DisplayMeshCache A8130A3E-E4F3-4CB0-BB8A-F10A473912D0    ON_BrepVertex[%d]:  ON_BrepEdge.m_brep = NULL (should point to parent ON_Brep)
 ON_BrepEdge.m_vi[1] = %d (should be >= 0 )
 ON_BrepEdge.m_vi[0] = %d (should be >= 0 )
 ON_BrepEdge.m_c3i = %d (should be >= 0 )
   ON_BrepEdge.m_edge_index = %d (should be >= 0 )
    ON_BrepEdge is not a valid curve proxy
 ON_BrepEdge[%d]:    trim.m_brep is null.
   trim.m_li = %d is not valid
    trim.m_iso = %d is not valid
   trim.m_type = ON_BrepTrim::slit is not valid. REserved for future use.
 trim.m_type = %d is not valid
  trim.m_v[1] = %d is not valid
  trim.m_v[0] = %d is not valid
  trim.m_ei = %d but trim.mtype != singular
  trim curve proxy settings are not valid.
   trim.m_c2i = %d is not valid
   trim.m_trim_index < 0.
 ON_BrepTrim[%d]:
   brep.m_L[%d] loop is not valid.
     )   (  ON_BrepFace[%d]:    ON_Brep.m_T[%d].m_pbox does not contain middle of trim.
    ON_Brep.m_T[%d].m_pbox does not contain end of trim.
   ON_Brep.m_T[%d].m_pbox does not contain start of trim.
 l�0=�#	@��0����� @�����`�D��2P2 ���0��`���� 	@	�	loop.m_type = %d is not a valid value.
 loop.m_brep is NULL.
   loop.m_fi = %d (should be >= 0 ).
  loop.m_ti[] is empty.
  loop.m_loop_index < 0.
 ON_BrepLoop[%d]: m_fi = %d, m_type = %d m_ti.Count() = %d
  ON_BrepFace m_brep = 0.  Should point to parent brep.
  ON_BrepFace m_si = %d.  Should be >= 0.
    ON_BrepFace m_li.Count() = 0  Should be > 0.
   ON_BrepFace m_face_index = %d.  Should be >= 0.
    ��<��<�    brep trim_index = %d (should be >=0 and <%d=brep.m_T.Count()).
 trim.m_c2i = %d (should be >=0 and <%d).
   trim.m_vi[0] = %d (should be >= 0 and < %d=brep.m_V.Count()).
  trim.m_vi[1] = %d (should be >= 0 and < %d=brep.m_V.Count()).
  trim.m_li = %d (should be >= 0 and <brep.m_L.Count()=%d
    trim.m_type = garbage (should be set to the correct ON_BrepTrim::TYPE value)
   trim.m_type = type_count (should be set to the correct ON_BrepTrim::TYPE value)
        trim.m_type = ON_BrepTrim::slit (should be set to the correct ON_BrepTrim::TYPE value)
 trim.m_brep does not point to parent brep.
 trim.m_pbox is not valid.
  trim.m_tolerance[1] = %g (should be >= 0.0)
    trim.m_tolerance[0] = %g (should be >= 0.0)
    trim.m_type = singular but trim.m_iso != N/S/E/W_iso
   trim.m_type = seam, the edge is manifold, but brep.m_L[trim.m_li=%d].m_type is not outer.
  edge.m_ti[%d]=%d is not a valid m_T[] index.
   All three trims have m_type = seam m_ei=%d and m_li = %d.
  brep.m_T[%d,%d, or %d] trim is not valid.
  edge.m_ti[%d] = m_ti[%d] = %d.
 brep.m_E[%d] trim is not valid.
    trim.m_type = seam but its other trim is not in the loop.
  trim.m_type = seam but brep.m_E[trim.m_ei=%d] < 2.
 trim.m_type = mated but brep.m_L[trim.m_li=%d].m_type is not inner or outer.
   trim.m_type = mated but brep.m_E[trim.m_ei=%d] only references this trim.
      trim.m_type = boundary but brep.m_L[trim.m_li=%d].m_type is not inner or outer.
        trim.m_type = boundary but brep.m_E[trim.m_ei=%d] has 2 or more trims.
 trim.m_type = unknown (should be set to the correct ON_BrepTrim::TYPE value)
   brep.m_E[trim.m_ei=%d].m_ti[] does not reference the trim.
     trim.m_type != singular and trim.m_ei = %d (m_ei should be >=0 and <brep.m_E.Count()=%d
        trim.m_type!=seam but brep.m_E[trim.m_ei=%d] references two trims in loop trim.m_li=%d.
    trim index %d is not in brep.m_E[trim.m_ei=%d].m_ti[]
      trim.m_vi[] = [%d,%d] but brep.m_C2[trim.m_c2i=%d]->IsClosed()=true
    trim.m_vi[1] != brep.m_E[trim.m_ei=%d].m_vi[trim.m_bRev3d?0:1]
 trim.m_vi[0] != brep.m_E[trim.m_ei=%d].m_vi[trim.m_bRev3d?1:0]
 trim.m_type = singular but brep.m_C2[trim.m_c2i=%d]->IsClosed() is true.
       trim.m_type = singular but trim.m_vi[] = [%d,%d] (the m_vi[] values should be equal).
  trim.m_type = singular but trim.m_ei = %d (should be -1)
       trim.Domain() = (%g,%g) is not included in brep.m_C2[trim.m_c2i=%d]->Domain() = (%g,%g)
    trim.Domain() = (%g,%g) (should be an increasing interval).
    trim.ProxyCurve() != m_C2[trim.m_c2i].
     trim.m_c2i = %d and ON_Brep.m_C2[%d]->Dimension() = %d (should be 2).
  trim.m_c2i = %d and ON_Brep.m_C2[%d] is NULL
   trim.m_trim_index = %d (should be %d).
 brep.m_T[%d] trim is not valid.
        brep loop_index = %d (should be >=0 and <%d=brep.m_L.Count()).
 loop.m_fi = %d (should be >= 0 and <brep.m_F.Count()=%d
    of brep.m_T[loop.m_ti[%d]=%d]=(%g,%g) do not match.
    end of brep.m_T[loop.m_ti[%d]=%d]=(%g,%g) and start 
       �����|�=loop.m_type = slit but loop has %d trims
       brep.m_T[loop.m_ti[%d]=%d].m_iso = E/W/N/S_iso (should be interior)
    brep.m_T[loop.m_ti[%d]=%d].m_type = %d (should be %d = seam)
   brep.m_L[%d] slit loop is not valid.
   brep.m_T[loop.m_ti[%d]=%d].m_li=%d (m_li should be %d).
    brep.m_T[loop.m_ti[%d]=%d] is not valid.
   loop.m_ti[%d] = loop.m_ti[%d] = %d (trim index can only appear once)
   loop.m_pbox is not valid
   loop.m_brep does not point to parent brep.
 loop.m_L[%d] loop is not valid.
    loop.m_type = %d (must be %d=outer, %d=inner, or %d=slit)
  loop.m_ti.Count() is <= 0  (should be > 0)
 loop.m_loop_index = %d (should be %d).
     brep face_index = %d (should be >=0 and <%d=brep.m_F.Count()).
 face.m_si=%d (should be >=0 and <%d=m_S.Count())
   face.ProxySurfaceIsTransposed() is true.
   brep.m_S[face.m_si=%d] != face.ProxySurface().
 brep.m_L[face.m_li[%d]=%d].m_type is not inner or slit.
    face.m_li[%d]=%d but brep.m_L[%d].m_fi=%d (m_fi should be %d)
  face.m_li[%d]=%d is a deleted loop
 brep.m_L[face.m_li[%d]=%d] is not valid.
       face.m_li[%d]=face.m_li[%d]=%d (a loop index should appear once in face.m_li[])
    brep.m_S[face.m_si=%d] is NULL
 brep.m_L[face.m_li[0]=%d].m_type is not outer.
 face.m_li.Count() <= 0 (should be >= 1)
    face.m_brep does not point to parent brep.
 face.m_face_index = %d (should be %d).
 brep.m_F[%d] face is not valid.
    brep edge_index = %d (should be >=0 and <%d=brep.m_E.Count() ).
    edge.m_c3i = %d (should be >=0 and <%d=m_C3.Count()
    edge.m_curve != brep.m_C3[edge.m_c3i=%d]
   edge.m_vi[0]=%d (should be >=0 and <%d=m_V.Count()
 edge.m_vi[1]=%d (should be >=0 and <%d=m_V.Count()
 edge.m_ti[%d]=%d (should be >=0 and <%d=m_T.Count())
   edge.m_ti[%d]=%d but brep.m_T[%d].m_ei=%d
      edge.m_ti[%d]=edge.m_ti[%d]=%d (a trim should be referenced once).
 edge.m_ti[%d]=%d is a deleted trim
 edge.m_tolerance=%g (should be >= 0.0)
 edge.m_ti.Count() < 0
  edge.m_vi[0]=edge.m_vi[1]=%d but edge.IsClosed() is false.
 edge.m_vi[%d]=%d but edge is not referenced in m_V[%d].m_ei[]
  edge.m_vi[%d]=%d is a deleted vertex
   edge.m_vi[]=(%d,%d) but edge.IsClosed() is true
    edge.m_domain=(%g,%g) is not valid
 edge is not a valid.
   edge.m_edge_index = %d (should be %d).
 edge.m_brep does not point to parent brep
  brep.m_E[%d] edge is not valid.
        brep vertex_index = %d (should be >=0 and <%d=brep.m_V.Count() ).
  vertex.m_ei[%d] = %d (should be >=0 and <%d).
      vertex.m_ei[%d] = %d but ON_Brep.m_E[%d].m_vi[] = [%d,%d]. At least one edge m_vi[] value should be %d.
        and ON_Brep.m_E[%d].m_vi[1] = %d (both m_vi[] values should be %d).
    vertex.m_ei[%d] and vertex.m_ei[%d] = %d but brep.m_E[%d].m_vi[0] = %d  in vertex.m_ei[] and a closed edge index should appear twice.
  vertex.m_ei[%d,%d,%d] = %d. An open edge index should appear once
  vertex.m_ei[%d] = %d is a deleted edge.
    vertex.m_tolerace = %g (should be >= 0.0)
  vertex.m_vertex_index = %d (should be %d).
 brep.m_V[%d] vertex is not valid.
  ON_Brep.m_T[%d] 2d curve is not inside surface domain.
 Bogus loop index in face.m_li[] .\opennurbs_brep.cpp    Bogus loop index in loop.m_ti[] Bogus trim.m_ei or trim.m_type value    Bogus loop index in trim.m_li   ON_Brep::IsManifold Bogus loop index in other_trim.m_li ON_Brep::LoopIsSurfaceBoundary  Bogus trim index in loop.m_ti[] ON_BrepEdge::EdgeCurveOf    ON_BrepEdge ProxyCurve() is NULL but m_c3i is valid ON_BrepTrim::TrimCurveOf    ON_BrepTrim ProxyCurve() = NULL but m_c2i is valid  d��V`V`�����p�0� � �W���	@�p���� � ��8 r@�0/0/��W��qON_BrepVertex m_ei[%d] = %d.  m_ei[] values should be >= 0
 ON_BrepVertex m_vertex_index = %d.  Should be >= 0
 <�`���� ����`
�Щ�p��@�!�P]@��
�
�n�W��0p 0 !	�<�=�. ��%p�>p��
�P� ��A�AP�@G� ���    ��0��� � �`�@����0�p����!�P]@��
�
�n�W�00p 0 !	�<�=�. ��%p�>p���P�@���AP�@G� ���    ,��� ��� PP �P����W���� r@��
�
�n�W�Pq|�p���� �@���P����W���!0B r����
�
�n���k�B!��!p"�" #�Y@#�#%$p&�#�&p' '�'�@�`(�( !	�B k )P)p)�)ON_Brep::AddTrimCurve   ON_Brep::AddTrimCurve() go a non-2d curve - changing dim to 2.  ON_Brep::AddEdgeCurve   ON_Brep::AddEdgeCurve() got a non-3d curve - changing dim to 3. ON_Brep.m_T[%d] is a seam trim with no matching seam trim in the same loop.
    Seam trim ON_Brep.m_T[%d].m_iso = W_iso but matching seam ON_Brep.m_T[%d].m_iso != E_iso.
      ON_Brep.m_T[%d,%d,%d] are three seam trims with the same edge in the same loop.
    ON_Brep.m_T[%d] is a seam trim with an invalid m_ei.
       Seam trim ON_Brep.m_T[%d].m_iso = N_iso but matching seam ON_Brep.m_T[%d].m_iso != S_iso.
      Seam trim ON_Brep.m_T[%d].m_iso = E_iso but matching seam ON_Brep.m_T[%d].m_iso != W_iso.
      Seam trim ON_Brep.m_T[%d].m_iso = S_iso but matching seam ON_Brep.m_T[%d].m_iso != N_iso.
      ON_Brep.m_F[%d] is on a closed surface. Outer loop m_L[%d] contains boundary trims %d and %d.  They should be seam trims connected to the same edge.
   ON_Brep.m_L[%d].m_pbox does not contain m_T[loop.m_ti[%d]].m_pbox.
     ON_Brep.m_L[%d] loop has trim vertex mismatch:
  m_T[loop.m_ti[%d]=%d].m_vi[1] = %d != m_T[loop.m_ti[%d]=%d].m_vi[0]=%d.
   ON_Brep.m_L[%d].m_pbox.m_max.z = %g (should be zero).
  ON_Brep.m_L[%d].m_pbox.m_min.z = %g (should be zero).
  ON_Brep.m_T[%d].m_vi[0] = %d is not invalid.
   ON_Brep.m_T[%d].m_vi[1] = %d is not invalid.
   ON_Brep.m_T[%d].m_c2i = %d is not valid.
   ON_Brep.m_T[%d].m_li = %d is not valid.
    ON_Brep.m_T[%d].m_ei = %d is not invalid.
  ON_Brep.m_T[%d].m_type = ON_BrepTrim::seam but m_iso is not N/E/W/S_iso.
   ON_Brep.m_T[%d].m_pbox.m_max.z = %g (should be zero).
  ON_Brep.m_T[%d].m_pbox.m_min.z = %g (should be zero).
      Distance from end of ON_Brep.m_T[%d] to 3d edge is %g.  (edge tol = %g, trim tol ~ %g).
        Distance from start of ON_Brep.m_T[%d] to 3d edge is %g.  (edge tol = %g, trim tol ~ %g).
      ON_Brep.m_T[%d].m_bRev3d = false, but closed curve directions are opposite.
    ON_Brep.m_T[%d].m_bRev3d = true, but closed curve directions are the same.
     ON_Brep.m_T[%d].m_bRev3d = %d, but m_vi[0] != m_E[m_ei].m_vi[%d].
  ON_Brep.m_T[%d].m_ei is deleted.
   ON_Brep.m_T[%d].m_iso = %d and it should be %d
 ON_Brep.m_T[%d].m_li = %d is a deleted loop.
   ON_Brep.m_T[%d].m_c2i = %d, but m_C2[%d] is NULL.
  ON_Brep.m_T[%d].m_vi[1] is deleted.
    ON_Brep.m_T[%d].m_vi[0] is deleted.
    ON_Brep.m_L[%d].m_fi = %d is not invalid.
  ON_Brep.m_L[%d].m_ti[%d] = %d is not invalid.
  ON_Brep.m_L[%d].m_ti[%d] = %d is a deleted trim.
   ON_Brep.m_L[%d].m_fi = %d is a deleted face.
   ON_Brep.m_F[%d] is invalid.
    ON_Brep.m_E[%d] is invalid.
    ON_Brep.m_V[%d] is invalid.
    ON_Brep.m_S[%d]->Dimension() = %d (should be 3).
   ON_Brep.m_S[%d] is invalid.
    ON_Brep.m_C3[%d] is a nested polycurve.
    ON_Brep.m_C3[%d]->Dimension() = %d (should be 3).
  ON_Brep.m_C3[%d] is invalid.
   ON_Brep.m_C2[%d] is a nested polycurve.
    ON_Brep.m_C2[%d]->Dimension() = %d (should be 2).
  ON_Brep.m_C2[%d] is invalid.
   ON_Brep.m_F[%d].m_face_index = %d (should be %d)
       ON_Brep.m_F[%d] is deleted (m_face_index = -1) but face.ProxySurface() is not NULL.
    ON_Brep.m_F[%d] is deleted (m_face_index = -1) but face.m_si=%d (should be -1).
        ON_Brep.m_T[%d].m_type = singular, but m_ei = %d (should be -1).
   ON_Brep.m_L[%d].m_loop_index = %d (should be %d)
   ON_Brep.m_L[%d] is deleted (m_loop_index = -1) but loop.m_fi=%d (should be -1).
        ON_Brep.m_F[%d] is deleted (m_face_index = -1) but face.m_li.Count()=%d.
   ON_Brep.m_T[%d] is not valid
   ON_Brep.m_T[%d].m_trim_index = %d (should be %d)
   ON_Brep.m_T[%d] is deleted (m_trim_index = -1) but trim.m_vi[0]=%d (should be -1).
     ON_Brep.m_T[%d] is deleted (m_trim_index = -1) but trim.m_c2i=%d (should be -1).
       ON_Brep.m_T[%d] is deleted (m_trim_index = -1) but trim.m_li=%d (should be -1).
        ON_Brep.m_T[%d] is deleted (m_trim_index = -1) but trim.m_ei=%d (should be -1).
        ON_Brep.m_L[%d] is deleted (m_loop_index = -1) but loop.m_ti.Count()=%d.
   ON_Brep.m_E[%d].m_edge_index = %d (should be %d)
   ON_Brep.m_E[%d] is deleted (m_edge_index = -1) but edge.m_vi[0]=%d (should be -1).
     ON_Brep.m_E[%d] is deleted (m_edge_index = -1) but edge.m_curve is not NULL.
   ON_Brep.m_E[%d] is deleted (m_edge_index = -1) but edge.m_c3i=%d (should be -1).
       ON_Brep.m_E[%d] is deleted (m_edge_index = -1) but edge.m_ti.Count() = %d.
     ON_Brep.m_T[%d] is deleted (m_trim_index = -1) but trim.m_vi[1]=%d (should be -1).
 ON_Brep.m_V[%d].m_vertex_index = %d (should be %d)
 ON_Brep.m_E[%d] is deleted (m_edge_index = -1) but edge.m_vi[1]=%d (should be -1).
     ON_Brep.m_V[%d] is deleted (m_vertex_index = -1) but vertex.m_ei.Count() = %d.
 ON_Brep has no vertices.
   ON_Brep has no 3d curves.
  ON_Brep has no 2d curves.
  ON_Brep has no trims.
  ON_Brep has no surfaces.
   ON_Brep has no loops.
  ON_Brep has no edges.
  ON_Brep has no faces, edges, or vertices
       j�t��?ON_Brep::CullUnusedSurfaces Brep face has illegal m_si. ON_Brep::CullUnused3dCurves Brep edge has illegal m_c3i.    ON_Brep::CullUnused2dCurves Brep trim has illegal m_c2i.    ON_Brep::CombineCoincidentVertices  ON_Brep::CombineCoincidentVertices - vertex0 = vertex1. domain(%g,%g) start(?,?) end(?,?)
  surface points start(%g,%g,%g) end(%g,%g,%g)
   domain(%g,%g) start(%g,%g) end(%g,%g)
  type(%s%s) rev3d(%d) 2d_curve(%d)
  trim[%2d]: edge(%2d) v0(%2d) v1(%2d) tolerance(%g,%g)
  -unknown_iso_flag   -north side iso -south side iso -v iso  -east side iso  -west side iso  -u iso  singular    seam        mated       boundary    unknown     loop[%2d]: type(%s) %d trims(   crvonsrf    slit    inner   outer   (Face geometry is the same as underlying surface.)
 Analysis mesh: %d polygons
 %s render mesh: %d polygons
    face[%2d]: surface(%d) reverse(%d) loops(   %s%d    ,%s%d   -   ?   trims ( domain(%g,%g) start(?,?,?) end(?,?,?)
  domain(%g,%g) start(%g,%g,%g) end(%g,%g,%g)
    edge[%2d]: v0(%2d) v1(%2d) 3d_curve(%d) tolerance(%g)
  edges ( vertex[%2d]: (%f %f %f) tolerance(%g)
  surface[%2d]: NULL
 surface details:
   surface[%2d]: %s u(%g,%g) v(%g,%g)
 curve3d[%2d]: %s domain(%g,%g) start(%g,%g,%g) end(%g,%g,%g)
   curve2d[%2d]: NULL
 curve2d[%2d]: %s domain(%g,%g) start(%g,%g) end(%g,%g)
 faces:     %d
  loops:     %d
  trims:     %d
  edges:     %d
  vertices:  %d
  2d curves: %d
  3d curve:  %d
  surfaces:  %d
  (B-rep geometry is the same as underlying surface.)
    ON_Brep:
   �����0�`�`� � �P� ���� �P� �h�����0�`��� � �P� ���������X�� �P� �����������`���@��fP�� � �����#��C r���]�
�
�E����p�B��L��@������Brep loop has illegal m_fi. ON_Brep::CullUnusedFaces    Brep face has illegal m_face_index. Brep trim has illegal m_li. Brep face m_li[] has illegal loop index.    ON_Brep::CullUnusedLoops    Brep loop has illegal m_loop_index. Brep edge.m_ti[] has illegal index. Brep loop.m_ti[] has illegal index. ON_Brep::CullUnusedTrims    Brep trim has illegal m_trim_index. Brep vertex.m_ei[] has illegal index.   Brep trim.m_ei has illegal index.   ON_Brep::CullUnusedEdges    Brep edge has illegal m_edge_index. Brep trim.m_vi[] has illegal index. Brep edge.m_vi[] has illegal index. Brep vertex has illegal m_vertex_index.     ON_Brep::CullUnusedVertices() - deleted vertex referenced by trim.m_vi[1]   ON_Brep::CullUnusedVertices ON_Brep::CullUnusedVertices() - deleted vertex referenced by trim.m_vi[0]   ON_BrepVertex   ON_Point    60B5DBC0-E660-11d3-BFE4-0010830122F0    ON_BrepEdge ON_CurveProxy   60B5DBC1-E660-11d3-BFE4-0010830122F0    ON_BrepTrim 60B5DBC2-E660-11d3-BFE4-0010830122F0    ON_BrepLoop 60B5DBC3-E660-11d3-BFE4-0010830122F0    ON_BrepFace ON_SurfaceProxy 60B5DBC4-E660-11d3-BFE4-0010830122F0    ON_Brep 60B5DBC5-E660-11d3-BFE4-0010830122F0    ON_Point::point is not a valid 3d point.
   ON_Point:   H��@ 0! ��`� 0��� � ��8 r@�0/0/��W��pqC3101A1D-F157-11d3-BFE7-0010830122F0    \������" ����`�0����� � �P� r@0��
�
�n�W��pq-- Attempting to continue.
 ERROR: Corrupt %s. (CRC errors).
   IDef    IDef_%02d   Layer   Layer_%02d  .\opennurbs_extensions.cpp  ��P�@(�(�(��a��<�<�p��( )�{����`)�)�)��`a��<���� *@*`/\�Pl ����(�� ��-.P.��`��. /@/4�0� *@*`/|����/0P0��Єp0 ��0� � 1`1�1T� �2P2 ���0��2 3����P�2P2 �,��`���8�7ONX_Model::Write archive.Write3dmEndMark() failed.
 ONX_Model::Write archive.EndWrite3dmHistoryTable() failed.
 ONX_Model::Write archive.BeginWrite3dmHistoryRecordTable() failed.
 ONX_Model::Write archive.EndWrite3dmObjectTable() failed.
  ONX_Model::Write archive.Write3dmObject(m_IDef_table[%d]) failed.
  ONX_Model::Write archive.BeginWrite3dmObjectTable() failed.
        ONX_Model::Write archive.EndWrite3dmInstanceDefinitionTable() failed.
  ONX_Model::Write archive.Write3dmInstanceDefinition(m_IDef_table[%d]) failed.
  ONX_Model::Write archive.BeginWrite3dmInstanceDefinitionTable() failed.
        ONX_Model::Write archive.EndWrite3dmHatchPatternTable() failed.
        ONX_Model::Write archive.Write3dmHatchPattern(m_hatch_pattern_table[%d]) failed.
       ONX_Model::Write archive.BeginWrite3dmHatchPatternTable() failed.
  ONX_Model::Write archive.EndWrite3dmLightTable() failed.
   ONX_Model::Write archive.Write3dmLight(m_light_table[%d]) failed.
  ONX_Model::Write archive.BeginWrite3dmLightTable() failed.
 ONX_Model::Write archive.EndWrite3dmDimStyleTable() failed.
    ONX_Model::Write archive.Write3dmDimStyle(m_dimstyle_table[%d]) failed.
    ONX_Model::Write archive.BeginWrite3dmDimStyleTable() failed.
  ONX_Model::Write archive.EndWrite3dmFontTable() failed.
    ONX_Model::Write archive.Write3dmFont(m_font_table[%d]) failed.
    ONX_Model::Write archive.BeginWrite3dmFontTable() failed.
  ONX_Model::Write archive.EndWrite3dmGroupTable() failed.
       ONX_Model::Write archive.Write3dmGroup(m_group_table[%d]) failed.
  ONX_Model::Write archive.BeginWrite3dmGroupTable() failed.
 ONX_Model::Write archive.EndWrite3dmLayerTable() failed.
       ONX_Model::Write archive.Write3dmLayer(m_layer_table[%d]) failed.
  ONX_Model::Write archive.BeginWrite3dmLayerTable() failed.
 ONX_Model::Write archive.EndWrite3dmLinetypeTable() failed.
    ONX_Model::Write archive.Write3dmLinetype(m_linetype_table[%d]) failed.
    ONX_Model::Write archive.BeginWrite3dmLinetypeTable() failed.
  ONX_Model::Write archive.EndWrite3dmMaterialTable() failed.
        ONX_Model::Write archive.Write3dmMaterial(m_material_table[%d]) failed.
    ONX_Model::Write archive.BeginWrite3dmMaterialTable() failed.
      ONX_Model::Write archive.EndWrite3dmTextureMappingTable() failed.
      ONX_Model::Write archive.Write3dmTextureMapping(m_mapping_table[%d]) failed.
   ONX_Model::Write archive.BeginWrite3dmTextureMappingTable() failed.
    ONX_Model::Write archive.EndWrite3dmBitmapTable() failed.
      ONX_Model::Write archive.Write3dmBitmap(m_bitmap_table[%d]) failed.
    ONX_Model::Write archive.BeginWrite3dmBitmapTable() failed.
    ONX_Model::Write archive.Write3dmSettings() failed.
Your m_settings information is not valid or basic file writing failed.
     ONX_Model::Write archive.Write3dmProperties() failed.
Your m_properties information is not valid or basic file writing failed.
 ONX_Model::Write archive.Write3dmStartSection() failed.
Your archive is not properly initialized
(make sure you passed ON::write3dm to the constructor),
a file is locked, a disk is locked, or something along those lines.
   ONX_Model::Write archive.Mode() is not ON::write3dm.
See ONX_Model::Write example in the header file.
  ONX_Model::Write version parameter = %d; it must be 0, or >= 2 and <= %d, or a multiple of 10 >= 50 and <= %d.
 ONX_Model::Write Your model is not valid and will not be saved.
    Duplicate object ids in model   ONX_Model::ObjectIndex  Nil object ids in model Duplicate idef ids in model ONX_Model::IDefIndex    Nil idef ids in model   Repaired.
  m_mapping_table[%d].m_mapping_index == %d (should be %d)
   m_group_table[%d].m_group_index == %d (should be %d)
   m_font_table[%d].m_font_index == %d (should be %d)
 m_dimstyle_table[%d].m_dimstyle_index == %d (should be %d)
 m_hatch_pattern_table[%d].m_hatchpattern_index == %d (should be %d)
    m_material_index = %d is not valid. m_linetype_index = %d is not valid.  Repaired.  m_layer_index = %d is not valid.    m_light_table[%d].m_attributes  m_light_table[%d].m_light_index == %d (should be %d)
   m_material_table[%d].MaterialIndex() == %d (should be %d)
  m_linetype_table[%d].LinetypeIndex() == %d (should be %d)
  m_layer_table[%d] and m_layer_table[%d] have same layer name.
  m_layer_table[%d].LayerName() is not valid
 m_layer_table[%d].LayerName() is empty
 m_layer_table[%d].LayerIndex() == %d (should be %d)
    m_idef_table[%d].m_object_uuid.Count() = 0.
    m_idef_table[%d].m_object_uuid[%d] is a circular reference.
        Object with uuid m_idef_table[%d].m_object_uuid[%d] has NULL m_object.
 Object with uuid m_idef_table[%d].m_object_uuid[%d] does not have m_attributes.Mode()=ON::idef_object.
 m_idef_table[%d].m_object_uuid[%d] is not an object's uuid.
    m_idef_table[%d].Name() = m_idef_table[%d].Name().
 m_idef_table[%d].Name() = "%ls" is not valid.
  m_object_table[%d].m_attributes m_object_table[%d].m_object->IsValid() = false.
    m_object_table[%d].m_object is NULL.
   t��l��<�wb  m_object_table[%d].m_attributes.m_uuid is nil.  m_object_table[%d] and [%d] have the same id.   m_light_table[%d] and m_object_table[%d] have same id.  m_light_table[%d] light id is nil.  m_light_table[%d] and[%d] have the same id. m_light_table[%d] light id and attributes id differ.    m_idef_table[%d].m_attributes.m_uuid is nil.    m_idef_table[%d] and[%d] are the same.  m_mapping_table[%d].m_mapping_id is nil.    m_mapping_table[%d] and[%d] are the same.   m_material_table[%d].m_material_id is nil.  m_material_table[%d] and[%d] are the same.  ��P� }p}�|�����0�p�T���`�Ђ��� �@�������`����� �8� � ������� ���������0�P�����P�������h� ����}�D@I G ' ��I`'D e f a u l t   ERROR: ON_BinaryArchive::Read3dmEndMark(&m_file_length) returned false.
        ERROR: Corrupt user data table. (ON_BinaryArchive::EndRead3dmUserTable() returned false.)
      ERROR: User data table entry %d is corrupt. (ON_BinaryArchive::Read3dmAnonymousUserTable() is false.)
  WARNING: Missing or corrupt history record table. (ON_BinaryArchive::BeginRead3dmHistoryRecordTable() returned false.)
 history record table    WARNING: Skipping history record table entry %d for unknown reason.
    ERROR: History record table entry %d is corrupt. (CRC errors).
 ERROR: History record table entry %d is corrupt. (ON_BinaryArchive::Read3dmHistoryRecord() < 0.)
       WARNING: Missing or corrupt object table. (ON_BinaryArchive::BeginRead3dmObjectTable() returned false.)
    object table        ERROR: Corrupt object light table. (ON_BinaryArchive::EndRead3dmObjectTable() returned false.)
 WARNING: Skipping object table entry %d for unknown reason.
    WARNING: Skipping object table entry %d because it's newer than this code.  Update your OpenNURBS toolkit.
     WARNING: Skipping object table entry %d because it's filtered.
 ERROR: Object table entry %d is corrupt. (CRC errors).
 ERROR: Object table entry %d is corrupt. (ON_BinaryArchive::Read3dmObject() < 0.)
      WARNING: Missing or corrupt instance definition table. (ON_BinaryArchive::BeginRead3dmInstanceDefinitionTable() returned false.)
   instance definition table   ERROR: Corrupt instance definition table. (ON_BinaryArchive::EndRead3dmInstanceDefinitionTable() returned false.)
      ERROR: Corrupt instance definition found. (ON_BinaryArchive::Read3dmInstanceDefinition() < 0.)
 WARNING: Missing or corrupt hatchpattern table. (ON_BinaryArchive::BeginRead3dmHatchPatternTable() returned false.)
    hatchpattern table      ERROR: Corrupt hatchpattern table. (ON_BinaryArchive::EndRead3dmHatchPatternTable() returned false.)
   ERROR: Corrupt hatchpattern found. (ON_BinaryArchive::Read3dmHatchPattern() < 0.)
      WARNING: Missing or corrupt render light table. (ON_BinaryArchive::BeginRead3dmLightTable() returned false.)
   render light table      ERROR: Corrupt render light table. (ON_BinaryArchive::EndRead3dmLightTable() returned false.)
  ERROR: Corrupt render light found. (ON_BinaryArchive::Read3dmLight() < 0.)
     WARNING: Missing or corrupt dimstyle table. (ON_BinaryArchive::BeginRead3dmDimStyleTable() returned false.)
    dimstyle table  ERROR: Corrupt dimstyle table. (ON_BinaryArchive::EndRead3dmDimStyleTable() returned false.)
   ERROR: Corrupt dimstyle found. (ON_BinaryArchive::Read3dmDimStyle() < 0.)
      WARNING: Missing or corrupt font table. (ON_BinaryArchive::BeginRead3dmFontTable() returned false.)
    font table      ERROR: Corrupt font table. (ON_BinaryArchive::EndRead3dmFontTable() returned false.)
   ERROR: Corrupt font found. (ON_BinaryArchive::Read3dmFont() < 0.)
      WARNING: Missing or corrupt group table. (ON_BinaryArchive::BeginRead3dmGroupTable() returned false.)
  group table     ERROR: Corrupt group table. (ON_BinaryArchive::EndRead3dmGroupTable() returned false.)
 ERROR: Corrupt group found. (ON_BinaryArchive::Read3dmGroup() < 0.)
    WARNING: Missing or corrupt layer table. (ON_BinaryArchive::BeginRead3dmLayerTable() returned false.)
  layer table     ERROR: Corrupt render layer table. (ON_BinaryArchive::EndRead3dmLayerTable() returned false.)
  ERROR: Corrupt layer found. (ON_BinaryArchive::Read3dmLayer() < 0.)
    WARNING: Missing or corrupt render linetype table. (ON_BinaryArchive::BeginRead3dmLinetypeTable() returned false.)
 render linetype table       ERROR: Corrupt render linetype table. (ON_BinaryArchive::EndRead3dmLinetypeTable() returned false.)
    ERROR: Corrupt render linetype found. (ON_BinaryArchive::Read3dmLinetype() < 0.)
       WARNING: Missing or corrupt render material table. (ON_BinaryArchive::BeginRead3dmMaterialTable() returned false.)
 render material table       ERROR: Corrupt render material table. (ON_BinaryArchive::EndRead3dmMaterialTable() returned false.)
    ERROR: Corrupt render material found. (ON_BinaryArchive::Read3dmMaterial() < 0.)
       WARNING: Missing or corrupt render texture_mapping table. (ON_BinaryArchive::BeginRead3dmTextureMappingTable() returned false.)
    render texture_mapping table        ERROR: Corrupt render texture_mapping table. (ON_BinaryArchive::EndRead3dmTextureMappingTable() returned false.)
       ERROR: Corrupt render texture_mapping found. (ON_BinaryArchive::Read3dmTextureMapping() < 0.)
  WARNING: Missing or corrupt bitmap table. (ON_BinaryArchive::BeginRead3dmBitmapTable() returned false.)
    bitmap table        ERROR: Corrupt bitmap table. (ON_BinaryArchive::EndRead3dmBitmapTable() returned false.)
       ERROR: Corrupt bitmap found. (ON_BinaryArchive::Read3dmBitmap() < 0.)
  settings section        ERROR: Unable to read settings section. (ON_BinaryArchive::Read3dmSettings() returned false.)
  properties section      ERROR: Unable to read properties section. (ON_BinaryArchive::Read3dmProperties() returned false.)
  start section       ERROR: Unable to read start section. (ON_BinaryArchive::Read3dmStartSection() returned false.)
      �V@��cܥL@��{��Ϊ?.\opennurbs_light.cpp   ON_Light::IsValid   ON_Light::IsValid(): illegal light style.   spot angle = %g degrees
    specular rgb =  diffuse rgb =   ambient rgb =   intensity = %g%%
   width =     length =    direction =     location =  index = %d  style = %s
 ambient_light   rectangular_light   linear_light    world_spot_light    world_point_light   world_directional_light camera_spot_light   camera_point_light  camera_directional_light              �?      (@ON_Light    85A08513-F383-11d3-BFE7-0010830122F0        �;f���?}Ô%�I�T��p��0P# �� �0��P�p#�W� �ON_Texture m_type has invalid value.
   ����1 ' ` 	���Ё�W  �@�ON_TextureMapping m_texture_space = %d is not a valid value.
   ON_TextureMapping m_projection = %d is not a valid value.
  ON_TextureMapping m_type = %d is not a valid value.
    UVW transformation:
    XYZ normal transformation:
 XYZ point transformation:
  single texture space
   divided texture space
  texture_space:  no projection
  closest point to mesh vertex
   mesh normal ray intersection
   projection:     %d
 box mapping
    sphere mapping
 cylinder mapping
   plane mapping
  no mapping
 type:   Texture mapping id:          �      ��      @    �?      @H��6�0ptexture[%d]:
   plug-in id =    index of refraction = %g
   reflectivity = %g%%
    transparency = %g%%
    shine = %g%%
   transparent rgb =   reflection rgb =    emmisive rgb =  id =    ON_RenderingAttributes error: m_materials[%d] and m_materials[%d] have the same plug-in id.
    ON_ObjectRenderingAttributes error: m_mappings[%d] and m_mappings[%d] have the same plug-in id.
    ���6P8�8�7��@��=p> �r�`� 4�E`�  �ON_Material 60B5DBBC-E660-11d3-BFE4-0010830122F0    ON_Texture  D6FF106D-329B-4f29-97E2-FD282A618020    ON_TextureMapping   32EC997A-C3BF-4ae5-AB19-FD572B8AD554    .\opennurbs_wstring.cpp w2c_size    Wide char string is not valid.  w2c     Error converting UTF-16 encoded wchar_t string to UTF-8 encoded char string.    c2w     Error converting UTF-8 encoded char string to UTF-16 encoded wchar_t string.    ON_wString::Empty   ON_wString::Empty() encountered invalid header - fixed.   	 
       {�G�zt?     @�@-C��6?-C��6?      4@      4�(��[�t`u @b��`�`z�u�W� � ��� r@���
�
�n�W��pqinvalid viewport port extents settings.
    invalid viewport frustum settings.
 invalid viewport camera settings.
  ON_Viewport::SetFrustum - invalid input .\opennurbs_viewport.cpp    ON_Viewport::SetFrustum ON_Viewport::SetFrustum - Beyond float precision perspective frus_near/frus_far values - will crash MS OpenGL      @ ؗA�G�z��?ON_Viewport.m_bValidFrustum in file was true and it should be false.    ON_Viewport::Read       ON_Viewport.m_bValidCamera in file was true and it should be false.           �?far: %d
    near: %d
   top: %d
    bottom: %d
 right: %d
  left: %d
   Port: (m_bValidPort = %s
   suggested minimum near/far: = %g
   suggested minimum near: = %g
   near/far: %g
   aspect (width/height):  far:    near:   top:    bottom:     right:  left:   top/bottom symmetry locked = %s
    left/right symmetry locked = %s
    Frustum: (m_bValidFrustum = %s)
    target distance %g
 Target Point:   Z:  Y:  X:  Direction:  (locked)    Camera: (m_bValidCamera = %s)
  parallel
   perspective
    invalid
    Projection:     ON_Viewport
    ON_Viewport D66E5CCF-EA39-11d3-BFE5-0010830122F0        �LX�z�ۿUnit system: %ls
   unknown unit system user defined unit (= %g meters) %ls (= %g meters)   parsecs light years astronomical units  nautical miles  picas (1/6 inch)    points (1/72 inch)  miles   yards   feet    inches  mils (= 0.001 inches)   microinches gigameters  megameters  kilometers  hectometers dekameters  meters  centimeters decimeters  millimeters microns nanometers  angstroms   no units    .\opennurbs_3dm_settings.cpp    ON_3dmUnitsAndTolerances::Write     ON_3dmUnitsAndTolerances::Write() - m_distance_display_precision out of range.        R@ON_3dmView::TargetPoint Obsolete ON_3dmView::m_target is not set correctly      �������x�P��� �����@����P����p�����P����P���relative viewport window position in application frame window
  left   = %6.2f%%, right = %6.2f%%
  bottom = %6.2f%%, top   = %6.2f%%
  viewport window screen location
  left   = %4d, right = %4d
  bottom = %4d, top   = %4d
  near   = %4d, far   = %4d
    view frustum
  left   = %g, right = %g
  bottom = %g, top   = %g
  near   = %g, far   = %g
 camera target
  distance = %g
  point = %g,%g,%g
   viewport camera frame
  location = %g, %g, %g
  X = %g, %g, %g
  Y = %g, %g, %g
  Z = %g, %g, %g
   Viewport: name = "%ls" projection = %s
 parallel    perspective     ON_3dmSettings::Read_v2() - TCODE_SETTINGS_CURRENT_FONT_INDEX - invalid font index value        ON_3dmSettings::Read_v2() - TCODE_SETTINGS_CURRENT_DIMSTYLE_INDEX - invalid dimstyle index value        ON_3dmSettings::Read_v2() - TCODE_SETTINGS_CURRENT_WIRE_DENSITY - invalid current_wire_density value    ON_3dmSettings::Read_v2 ON_3dmSettings::Read_v2() - TCODE_SETTINGS_CURRENT_LAYER_INDEX - invalid layer index value  ��0	� 	 ������	�#	@��0(�p	0��:0�t��	�� �  � ��@� ����(��		`V`���X���`V`������		0��:0���
	���8�7t��	�#	@��0.\opennurbs_archive.cpp DownSizeINT i64 too big to convert to 4 byte signed int DownSizeUINT    u64 too big to convert to 4 byte unsigned int       ��0	 1	02	 @��0����i	�W� �p	�W�OBSOLETE CustomMeshUserData ON_BinaryArchive::SetArchive3dmVersion  ON_BinaryArchive::SetArchive3dmVersion - invalid version    ON_BinaryFile::CurrentPosition() NULL file. ON_BinaryFile::CurrentPosition  ON_BinaryFile::CurrentPosition() - _ftelli64() failed   ON_BinaryFile::SeekFromCurrentPosition  ON_BinaryFile::Seek() fseek(,SEEK_CUR) failed.  ON_BinaryFile::SeekFromStart    ON_BinaryFile::SeekFromStart() fseek(,SEEK_SET) failed. ,�0%	�#	@��0�Z�1�q�I�uuu��7�ON_BinaryArchive::FindMisplacedTable        ON_BinaryArchive::FindMisplacedTable - must provide plug-in id when searching for user tables   ON_BinaryArchive::ReadByte() NULL file or buffer.   ON_BinaryArchive::ReadByte() Read() failed. ON_BinaryArchive::ReadByte  ON_BinaryArchive::ReadByte() ReadMode() is false.   ON_BinaryArchive::WriteByte() NULL file or buffer.  ON_BinaryArchive::WriteByte() fwrite() failed.  ON_BinaryArchive::WriteByte ON_BinaryArchive::WriteByte() WriteMode() is false. t��p	���������������]
ON_BinaryArchive::ReadTime  ON_BinaryArchive::ReadTime() - bad time in archive  string element count is impossibly large    string byte count exceeds current chunk size    ON_BinaryArchive::ReadStringUTF16ElementCount   ON_BinaryArchive::ReadBool  ON_BinaryArchive::ReadBool - bool value != 0 and != 1       ON_BinaryArchive::EndRead3dmChunk: partially read chunk - skipping bytes at end of current chunk.       ON_BinaryArchive::EndRead3dmChunk: current position after end of current chunk. ON_BinaryArchive::EndRead3dmChunk: CRC32 error. ON_BinaryArchive::EndRead3dmChunk: current position before start of current chunk.  ON_BinaryArchive::EndRead3dmChunk: CRC16 error. ON_BinaryArchive::EndRead3dmChunk   ON_BinaryArchive::EndRead3dmChunk - negative chunk length   ON_BinaryArchive::Read3dmAnonymousUserTable ON_BinaryArchive::Read3dmAnonymousUserTable() do not read a TCODE_USER_RECORD chunk.    �� �	�	�	P	P	`	�	@	�]
� �	 	  	` 	� 	� 	 !	�
�]
ON_BinaryArchive::EndWrite3dmChunk() - CurrentPosition() != offset  ON_BinaryArchive::EndWrite3dmChunk() - chunk length < 0 ON_BinaryArchive::EndWrite3dmChunk  ON_BinaryArchive::EndWrite3dmChunk: CRC16 computation error.    ON_BinaryArchive::EndRead3dmTable() m_chunk.Last()->typecode != typecode        ON_BinaryArchive::EndRead3dmTable() v2 file m_chunk.Count() != 1        ON_BinaryArchive::EndRead3dmTable() v1 file m_chunk.Count() != 0    ON_BinaryArchive::EndRead3dmTable() m_active_table != t ON_BinaryArchive::EndRead3dmTable   ON_BinaryArchive::EndRead3dmTable() bad typecode    ON_BinaryArchive::EndRead3dmLayerTable() - m_chunk.Count() > 0  ON_BinaryArchive::EndRead3dmLayerTable      ON_BinaryArchive::EndRead3dmLayerTable() - m_active_table != no_active_table    ON_BinaryArchive::BeginRead3dmChunk() - file is damaged.    ON_BinaryArchive::BeginRead3dmBigChunk      ON_BinaryArchive::BeginRead3dmChunk() - Rogue eof marker in v2 file.
   ON_BinaryArchive::BeginRead3dmChunk - unexpected tcode or chunk length - archive driver or device may be bad    ON_BinaryArchive::BeginRead3dmChunk - minor_version < 0 ON_BinaryArchive::BeginRead3dmChunk - major_version < 1 ON_BinaryArchive::BeginRead3dmChunk - unexpected chunk length   ON_BinaryArchive::BeginRead3dmChunk - unexpected tcode  ON_BinaryArchive::BeginRead3dmChunk - input minor_version NULL  ON_BinaryArchive::BeginRead3dmChunk - input major_version NULL  ON_BinaryArchive::BeginRead3dmChunk - input expected_tcode has short flag set.  ON_BinaryArchive::BeginRead3dmChunk ON_BinaryArchive::BeginRead3dmChunk - input expected_tcode = 0  May 18 2015  (compiled on    3DM I/O processor: OpenNURBS toolkit version %d    3D Geometry File Format %8d 3dm archive version must be 2, 3, 4 or 50   ON_BinaryArchive::Write3dmStartSection      3dm archive version must be <= ON_BinaryArchive::CurrentArchiveVersion()        ON_BinaryArchive::Read3dmStartSection(): Archive has V1 header and V2 body. Continuing to read V2 body. ON_BinaryArchive::Read3dmStartSection   ON_BinaryArchive::Read3dmStartSection - start section string is unreasonably long.  3D Geometry File Format     http://www.rhino3d.com  Rhinoceros  Interface:  ON_BinaryArchive::Read3dmProperties Comment length > 1000000    ON_BinaryArchive::Read3dmV1Layer    ON_BinaryArchive::Read3dmV1Layer() - invalid layer name length  RhAnnotateDot   RhAnnotateArrow RhFreezePrevLayer   RhHidePrevLayer       P@ON_BinaryArchive::Read3dmV1Light    ON_BinaryArchive::Read3dmV1Light() m_chunk.Count() != 0          �_@    ���@ON_BinaryArchive::EndRead3dmTable() m_chunk.Last()->typecode != TCODE_USER_RECORD       ON_BinaryArchive::EndRead3dmTable() missing TCODE_ENDOFTABLE marker.    ON_BinaryArchive::EndRead3dmUserTable   ON_BinaryArchive::EndRead3dmUserTable() m_chunk.Count() != 2    Unable to read user data header information.    ReadObjectUserDataHeaderHelper  version 2.0 TCODE_OPENNURBS_CLASS_USERDATA chunk is missing TCODE_OPENNURBS_CLASS_USERDATA_HEADER chunk.        Unable to read TCODE_OPENNURBS_CLASS_USERDATA chunk version numbers Reading object user data - length of TCODE_ANONYMOUS_CHUNK < 4      Reading object user data - unable to find TCODE_ANONYMOUS_CHUNK Unable to create object user data class. Flawed class id information.   Reading object user data - unable to create userdata class  ON_BinaryArchive::ReadObjectUserData    TCODE_OPENNURBS_CLASS_USERDATA chunk is too short   ON_BinaryArchive::BeginWrite3dmChunk - input minor_version < 0. ON_BinaryArchive::BeginWrite3dmChunk - input major_version <= 0.        ON_BinaryArchive::BeginWrite3dmChunk - input tcode has short flag set.  ON_BinaryArchive::BeginWrite3dmChunk    ON_BinaryArchive::BeginWrite3dmChunk - input tcode = 0  ON_BinaryArchive::BeginWrite3dmTable() m_chunk.Count() > 0      ON_BinaryArchive::BeginWrite3dmTable() m_active_table != no_active_table    ON_BinaryArchive::BeginWrite3dmTable    ON_BinaryArchive::BeginWrite3dmTable() bad typecode ON_BinaryArchive::EndWrite3dmTable() m_chunk.Last()->typecode != typecode   ON_BinaryArchive::EndWrite3dmTable() m_chunk.Count() != 1   ON_BinaryArchive::EndWrite3dmTable() m_active_table != t    ON_BinaryArchive::EndWrite3dmTable  ON_BinaryArchive::EndWrite3dmTable() bad typecode       ON_BinaryArchive::BeginWrite3dmLayerTable() - m_active_table != no_active_table ON_BinaryArchive::BeginWrite3dmLayerTable       ON_BinaryArchive::BeginWrite3dmLayerTable() - chunk stack should be empty   ON_BinaryArchive::EndWrite3dmLayerTable     ON_BinaryArchive::EndWrite3dmLayerTable() - m_active_table != layer_table       ON_BinaryArchive::BeginWrite3dmUserTable() - nil usertable_uuid not permitted.  ON_BinaryArchive::BeginWrite3dmUserTable        ON_BinaryArchive::BeginWrite3dmUserTable() - m_active_table != no_active_table  ON_BinaryArchive::EndWrite3dmUserTable  ON_BinaryArchive::EndWrite3dmUserTable() - not in a TCODE_USER_RECORD chunk.    ON_BinaryArchive::Write3dmEndMark       ON_BinaryArchive::WriteEndMark() called with unfinished chunks.
        ON_UnknownUserData::Cast(ud) is not null and ud->IsUnknownUserData() is false.  ON_BinaryArchive::WriteObjectUserData   ON_UnknownUserData::Cast(ud) is null and ud->IsUnknownUserData() is true.   Not saving %s userdata - m_application_uuid is nil. ON_BinaryArchive::ReadObject() pObject->Read() failed.  ON_BinaryArchive::ReadObject() pID->Create() returned NULL.     ON_BinaryArchive::ReadObject() TCODE_OPENNURBS_CLASS_DATA chunk length too small        ON_BinaryArchive::ReadObject() didn't find TCODE_OPENNURBS_CLASS_DATA block     ON_BinaryArchive::ReadObject() ON_ClassId::ClassId(uuid) returned NULL. ON_BinaryArchive::ReadObject() - uuid does not match intput pObject's class id. ON_BinaryArchive::ReadObject() TCODE_OPENNURBS_CLASS_UUID has invalid length    ON_BinaryArchive::ReadObject() didn't find TCODE_OPENNURBS_CLASS_UUID block     ON_BinaryArchive::ReadObject() TCODE_OPENNURBS_CLASS chunk length too small.    ON_BinaryArchive::ReadObjectHelper      ON_BinaryArchive::ReadObject() didn't find TCODE_OPENNURBS_CLASS block. ON_BinaryArchive::Seek3dmChunkFromStart() called with out of bounds current position    ON_BinaryArchive::Seek3dmChunkFromStart() called with an active chunk that has m_value < 0  ON_BinaryArchive::Seek3dmChunkFromStart     ON_BinaryArchive::Seek3dmChunkFromStart() - current chunk is not a long chunk   ON_BinaryArchive::BeginRead3dmTable() - corrupt table - skipping        ON_BinaryArchive::BeginRead3dmTable() - current file position not at start of table - searching ON_BinaryArchive::BeginRead3dmTable() m_chunk.Count() > 0       ON_BinaryArchive::BeginRead3dmTable() m_active_table != no_active_table ON_BinaryArchive::BeginRead3dmTable ON_BinaryArchive::BeginRead3dmTable() bad typecode  ON_BinaryArchive::BeginRead3dmUserTable() - missing user table TCODE_USER_RECORD chunk. ON_BinaryArchive::BeginRead3dmUserTable ON_BinaryArchive::BeginRead3dmUserTable() - missing user table UUID ON_BinaryArchive::WriteObject() o.Write() failed.   ON_BinaryArchive::WriteObject   ON_BinaryArchive::WriteObject() o.ClassId() returned NULL.  ON_BinaryArchive::ReadObject    ON_BinaryArchive::ReadObject() called with NULL ppObject.   ON_BinaryArchive::Write3dmBitmap        ON_BinaryArchive::Write3dmBitmap() must be called in BeginWrite3dmBitmapTable() block   ON_BinaryArchive::Read3dmBitmap ON_BinaryArchive::Read3dmBitmap() - corrupt bitmap table        ON_BinaryArchive::Write3dmLayer() must be called in BeginWrite3dmLayerTable(2) block    ON_BinaryArchive::Write3dmLayer() - version 1 - chunk stack should be empty ON_BinaryArchive::Write3dmLayer     ON_BinaryArchive::Write3dmLayer() - m_active_table != layer_table   ON_BinaryArchive::Read3dmLayer() - corrupt layer table  ON_BinaryArchive::Read3dmLayer      ON_BinaryArchive::BeginRead3dmLayerTable() - m_active_table != no_active_table  ON_BinaryArchive::Write3dmGroup() must be called in BeginWrite3dmGroupTable() block ON_BinaryArchive::Write3dmGroup     ON_BinaryArchive::Write3dmGroup() - m_active_table != group_table   ON_BinaryArchive::Read3dmGroup() - corrupt group table  ON_BinaryArchive::Read3dmGroup      ON_BinaryArchive::BeginRead3dmGroupTable() - m_active_table != no_active_table  ON_BinaryArchive::Write3dmFont() must be called in BeginWrite3dmFontTable() block   ON_BinaryArchive::Write3dmFont      ON_BinaryArchive::Write3dmFont() - m_active_table != font_table ON_BinaryArchive::Read3dmFont() - corrupt font table    ON_BinaryArchive::Read3dmFont   ON_BinaryArchive::BeginRead3dmFontTable() - m_active_table != no_active_table   ON_BinaryArchive::Write3dmDimStyle() must be called in BeginWrite3dmDimStyleTable() block   ON_BinaryArchive::Write3dmDimStyle  ON_BinaryArchive::Write3dmDimStyle() - m_active_table != dimstyle_table ON_BinaryArchive::Read3dmDimStyle() - corrupt dimstyle table    ON_BinaryArchive::Read3dmDimStyle       ON_BinaryArchive::BeginRead3dmDimStyleTable() - m_active_table != no_active_table       ON_BinaryArchive::Write3dmHatchPattern() must be called in BeginWrite3dmHatchPatternTable() block   ON_BinaryArchive::Write3dmHatchPattern      ON_BinaryArchive::Write3dmHatchPattern() - m_active_table != hatchpattern_table ON_BinaryArchive::Read3dmHatchPattern() - corrupt hatch pattern table   ON_BinaryArchive::Read3dmHatchPattern   ON_BinaryArchive::BeginRead3dmHatchPatternTable() - m_active_table != hatchpattern_table        ON_BinaryArchive::Write3dmLinetype() must be called in BeginWrite3dmLinetypeTable() block   ON_BinaryArchive::Write3dmLinetype  ON_BinaryArchive::Write3dmLinetype() - m_active_table != linetype_table ON_BinaryArchive::Read3dmLinetype() - corrupt linetype table    ON_BinaryArchive::Read3dmLinetype       ON_BinaryArchive::BeginRead3dmLinetypeTable() - m_active_table != linetype_table        ON_BinaryArchive::Write3dmInstanceDefinition() must be called in BeginWrite3dmInstanceDefinitionTable() block   ON_BinaryArchive::Write3dmInstanceDefinition    ON_BinaryArchive::Write3dmInstanceDefinition() - m_active_table != instance_definition_table    ON_BinaryArchive::Read3dmInstanceDefinition() - corrupt instance definition table   ON_BinaryArchive::Read3dmInstanceDefinition ON_BinaryArchive::BeginRead3dmInstanceDefinitionTable() - m_active_table != no_active_table     ON_BinaryArchive::Write3dmTextureMapping() - active chunk typecode != TCODE_TEXTURE_MAPPING_TABLE   ON_BinaryArchive::Write3dmTextureMapping    ON_BinaryArchive::Write3dmTextureMapping() - m_active_table != texture_mapping_table    ON_BinaryArchive::Read3dmTextureMapping ON_BinaryArchive::Read3dmTextureMapping() - corrupt texture_mapping table       ON_BinaryArchive::Write3dmHistoryRecord() - active chunk typecode != TCODE_HISTORYRECORD_TABLE  ON_BinaryArchive::Write3dmHistoryRecord ON_BinaryArchive::Write3dmHistoryRecord() - m_active_table != history_record_table  ON_BinaryArchive::Read3dmHistoryRecord      ON_BinaryArchive::Read3dmHistoryRecord() - corrupt history_record table ON_BinaryArchive::Write3dmMaterial() - active chunk typecode != TCODE_MATERIAL_TABLE    ON_BinaryArchive::Write3dmMaterial      ON_BinaryArchive::Write3dmMaterial() - m_active_table != material_table ON_BinaryArchive::Read3dmMaterial   ON_BinaryArchive::Read3dmMaterial() - corrupt material table        ON_BinaryArchive::Write3dmMaterial() - active chunk typecode != TCODE_LIGHT_TABLE   ON_BinaryArchive::Write3dmLight     ON_BinaryArchive::Write3dmLight() - m_active_table != light_table   ON_BinaryArchive::Read3dmLight() - corrupt light table  ON_BinaryArchive::Read3dmLight      ON_BinaryArchive::Read3dmLight() - m_active_table != light_table        ON_BinaryArchive::Write3dmObject() - active chunk typecode != TCODE_OBJECT_TABLE    ON_BinaryArchive::Write3dmObject    ON_BinaryArchive::Write3dmObject() - m_active_table != object_table ON_BinaryArchive::Read3dmObject() - corrupt object table    ON_BinaryArchive::Read3dmObject ON_BinaryArchive::Read3dmObject() - missing TCODE_OBJECT_RECORD_TYPE chunk. ON_OBSOLETE_CCustomMeshUserData 69F27695-3011-4FBA-82C1-E529F25B5FD9        �C�h[C`#��=�@C  �+]jAB     �@L7�A`%�@     ��@��)A�B?�0��(?�eu����>�q�q�?UUUUUU�?��x�v�=?$�E[>��t�i�0?����d?     ��@    ,9xA    wG�A�5��B��>�
F%u�?���̋��<��Jw�<��-f�=��g|�A?    e��A��K7�A�?R���Q@ffffff9@T��Z
�P
`P
	   ON_UNSET_VALUE  UnsetPoint  >   <   UnsetVector zero transformation
    identity transformation
    %08X-%04X-%04x-%02X%02X-%02X%02X%02X%02X%02X%02X    %08X-...(runtime value varies)  %d %d %d    ON_UNSET_COLOR  December    November    October September   August  July    June    May April   March   February    January Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday   = (    %c  %s[%2d] %c  %sNULL point list
  %sEMPTY point list
 %s[%2d] point   %5d  %23.17g  %4d  %10.4g
  %5d  %23.17g  %4d
  index                     value  mult       delta
  knot vector cv_count < order
   knot vector order < 2
  NULL knot vector
   %.17g   %g      PolylineCurve m_t.Count() = %d and PointCount() = %d (should be equal)
 PolylineCurve has %d points (should be >= 2)
   PolylineCurve m_t[%d]=%g should be less than m_t[%d]=(%g).
 PolylineCurve m_dim = %d (should be 2 or 3).
   PolylineCurve m_pline[] is not valid.
  , %g
     point[%2d] =  ON_PolylineCurve:  domain = [%g,%g]
        �� \
�
��
 �`
�a
�_
�_
�\
 ]
p�� �0\
0`
0�@@\
0/0/p\
�W��p0p���b
�c
Ѝ
�d
�]
@f
=���=�f
@g
�]
�>�g
�h
�]
�W`i
 p
 r
�r
`s
 t
�v
��
��
��
�]
 ^
 ^
ON_PolylineCurve    4ED7D4E6-E947-11d3-BFE5-0010830122F0          �<Name: %ls
  .\opennurbs_3dm_properties.cpp  ON_SetBinaryArchiveOpenNURBSVersion ON_SetBinaryArchiveOpenNURBSVersion - invalid opennurbs version ON_3dmProperties::Read  ON_3dmProperties::Read - TCODE_PROPERTIES_OPENNURBS_VERSION corrupt value       openNURBS ERROR # %d - Too many errors.  No more printed messages.  openNURBS ERROR # %d %s.%d  openNURBS ERROR # %d %s.%d %s():        openNURBS WARNING # %d - Too many warnings.  No more printed messages.  openNURBS WARNING # %d %s.%d    openNURBS WARNING # %d %s.%d %s():    CV[%2d]   Knot Vector %d ( %d knots )
    ON_NurbsSurface dim = %d is_rat = %d
        order = %d X %d cv_count = %d X %d
    ON_NurbsSurface.m_cv_stride[] = {%d,%d} is not valid.
      ON_NurbsSurface.m_cv_stride[%d]=%d is too small (should be >= %d).
 ON_NurbsSurface.m_knot[%d] is not a valid knot vector.
 ON_NurbsSurface.m_knot[i] is NULL.
 ON_NurbsSurface.m_cv_count[%d] = %d (should be >= m_order[%d]=%d).
 ON_NurbsSurface.m_order[i] = %d (should be >= 2).
  ON_NurbsSurface.m_cv is NULL.
  ON_NurbsSurface.m_dim = %d (should be > 0).
    .\opennurbs_nurbssurface.cpp    ����
��������8��
`�
0�
 ��
�
 �
��
��
��
�W� �p1@�
 r@`�
0/0/�
���k�p�B���
з
@�
��
��
�YP�
�
 ^�Z@�
 �
 �
��
��
 �
P�
��
�
 �
��
 �
��
��
�Wkk�
ON_NurbsSurface::TensorProduct() - tensor.DimensionB() > dimB   ON_NurbsSurface::TensorProduct  ON_NurbsSurface::TensorProduct() - tensor.DimensionA() > dimA   ON_NurbsSurface 4ED7D4DE-E947-11d3-BFE5-0010830122F0        ����
�� ��
��
��
�
P � �W���
�� r�� 0�n���k�p�B��`��P
�
�Y�
 ^�Z�P��Pp��� �`�@ON_SumSurface.m_curve[%d] is not valid.
    ON_SumSurface.m_curve[%d]->m_dim = %d (should be 3).
   ON_SumSurface.m_curve[%d] is NULL.
 ON_SumSurface.m_basepoint is not valid.
    m_curve[%d] = NULL
 m_curve[%d]:
   basepoint =     ���6����ON_SumSurface   C4CD5359-446D-4690-9FF5-29059732472B    ,�0"PQ@_  %�&�#$ (�(�W�@" �`_ r�P0*�
�
�n���k�p�B��K�K�L O�O�Y�P`J ^�Z I J�H�G�E�D0E�D@, :�>pAY�R�I�6`8ON_RevSurface.m_t = (%g,%g) (should be an increasing interval)
 ON_RevSurface.m_angle.Length() = %g (should be > ON_ZERO_TOLERANCE).
   ON_RevSurface.m_angle.Length() = %g (should be <= 2*pi radians).
       -HT�!@ON_RevSurface.m_angle = (%g,%g) (should be an increasing interval)
 ON_RevSurface.m_axis is not valid.
 ON_RevSurface.m_curve->Dimension()=%d (should be 3).
   ON_RevSurface.m_curve is not valid.
    ON_RevSurface.m_curve is NULL.
 Revolute: 
 Angle evaluation parameter interval: [%g,%g].
  Rotation angle: %g to %g radians.
  Axis:   Paramerization: (angle,curve)
  Paramerization: (curve,angle)
  ���6� � � 5-@T�!@�*�`�!	@�*�`�!�?ON_RevSurface.m_curve is not valid. .\opennurbs_revsurface.cpp  ON_RevSurface::GetNurbForm  ON_RevSurface.m_curve is 2-dimensional. ON_RevSurface   A16220D3-163B-11d4-8000-0010830122F0        ��{��Ϊ?�� e��@� `�0��} ~���p���}0�P���@���0����W��p�B@�� ��P�����=���=������>�����`�������� � �`���P��� �`� �Polycurve segment count = %d and dim = %d
  Polycurve end of segment[%d] != start of segment[%d] (distance=%g)
 Polycurve segment[%d] is closed (%d segments).
 Polycurve m_t[%d]=%g and m_t[%d]=%g (should be increasing)
 Polycurve segment[%d]->Dimension()=%d (should be %d).
  Polycurve segment[%d] is not valid.
    Polycurve segment[%d] is null.
 Polycurve segment count = %d and m_t.Count()=%d (should be segment count+1)
    null curve pointer
  invalid previous segment curve  invalid segment curve   gap = %.17g    Segment %d: (%g,%g) ON_PolyCurve segment count = %d
    .\opennurbs_polycurve.cpp   +�����?ON_PolyCurve::Read  ON_PolyCurve::Read() - non ON_Curve object in segment list
 ON_PolyCurve    4ED7D4E0-E947-11d3-BFE5-0010830122F0     �P��W � @��0�����W� ��r�W�user data saved in 3dm archive: %s
 no  yes user data copy count: %d
   user data uuid:     user data description: %ls
 n o n e     User Data:
     invalid userdata - classes derived from ON_UserData that get saved in 3dm archives must have a class id and name defined by ON_OBJECT_DECLARE/ON_OBJECT_IMPLEMENT.
     invalid userdata - m_userdata_uuid in use. Use guidgen to get a unique id.
 invalid userdata - m_userdata_uuid = nil
   4������� ��p������ ��W� ������    Unknown user data. (Definition of class was not available when object was read.)    Data size in 3dm archive: %d bytes
 unknown class uuid:     ������ �@�p��� !	�
�]
Value: %ls
 Key: %ls
   ��P���p� �r �`��`����W� �User text (%d entries)  %d entries
     ��` �  @� �p����� �W� �@����850324A7-050E-11d4-BFFA-0010830122F0    ON_UnknownUserData  850324A8-050E-11d4-BFFA-0010830122F0    ON_UserStringList   CE28DE29-F4C5-4faa-A50A-C3A6849B6329    ON_DocumentUserStringList   06F3218E-F5EC-4f6c-B74C-14583F0ED7BC    l��#�g`; @� �p$��$0%�W� � &���Userdata extension of ON_TextEntity �� &�h�< @� �p'��'0(�W� �)���Userdata extension of ON_Dimensions < >     ��1�W�X @� �p2��2�2�W� ��3���Userdata extension of ON_AngularDimension2  A r i a l   b o l d     \��*�?Pd �6 7`�`7�7�8� � ��8 r@�0/0/�n�W��pqON_TextDot m_point is not valid
    ON_TextDot "%ls" at         ���8�d`9 @��0�����W� �0:�W�Annotation Text Formula ON_Annotation2 - m_type = %d is not a valid enum value
 ON_Annotation2 - m_points[%d] is not valid.
    ON_Annotation2 - m_plane is not valid
      ON_LinearDimension2 - m_points[3].y = %g != %g = m_points[1].y
 ON_LinearDimension2 - m_points[3].x = %g != %g = m_points[2].x
 ON_LinearDimension2 - m_points[1].x = %g != %g = m_points[0].x (should be equal)
   ON_LinearDimension2 - m_points.Count() = %d (should be 5).
 ON_LinearDimension2 - invalid ON_Annotation2 base class.
       ON_LinearDimension2 - m_type !=  ON::dtDimLinear or ON::dtDimAligned.
  R    �>ON_RadialDimension2 - m_points.Count() = %d (should be 4 or 5)
 ON_RadialDimension2 - invalid ON_Annotation2 base class.
       ON_RadialDimension2 - m_type !=  ON::dtDimRadius or ON::dtDimDiameter
  ON_AngularDimension2 - bogus m_angle = %g
  ON_AngularDimension2 - bogus m_radius = %g
 ON_AngularDimension2 - angle dim m_points[3] = not on arc interior.
    ON_AngularDimension2 - m_radius = %g != %g = |m_point[3])|
     ON_AngularDimension2 - m_angle = %g != %g = (end angle - start angle)
  ON_AngularDimension2 - angle dim m_points[3] = center (should be on interior of arc).
  ON_AngularDimension2 - angle dim m_points[2] = center (should be on end ray).
  ON_AngularDimension2 - angle dim m_points[1] = center (should be on start ray).
    ON_AngularDimension2 - m_points.Count() = %d (should be 4)
 ON_AngularDimension2 - invalid ON_Annotation2 base class.
  ON_AngularDimension2 - m_type !=  ON::dtDimAngular
 ON_OrdinateDimension2 - m_points.Count() = %d (should be 2).
   ON_OrdinateDimension2 - invalid ON_Annotation2 base class.
 ON_OrdinateDimension2 - m_type !=  ON::dtDimOrdinate.
      �������?ON_Leader2 - m_points.Count() = %d (should be >= 2)
    ON_Leader2 - invalid ON_Annotation2 base class.
    ON_Leader2 - m_type !=  ON::dtLeader
       ��0)�W0� �@�`�P�pk �� � ��� r@���
�
�n�W��p�j`1pM�1�1L�p) �P� �M�`���} �� � � n�p@@S�
�
�n�W��p�j VpM�1�1���)� � @V�`���} �� � ��q t@P��
�
�n�W��p�j�VpM�1�1���) �`� �X�`���Pw �� � � upv@�A�
�
�n�W��p�j�3pM�1�1H�P+ �`� �`�`���x �� � � y�z@`��
�
�n�W��p�jpapM�1�1��0* �P�  |�`���} �� � ��a�}@�3�
�
�n�W��p�j`1pM�5�5ON_TextEntity2 - m_points.Count() = %d (should be 0)
   ON_TextEntity2 - invalid ON_Annotation2 base class.
    ON_TextEntity2 - m_usertext does not contain printable characters.
 ON_TextEntity2 - m_type !=  ON::dtTextBlock
        ��p* ��� �c�`���} �� � ��~`�@��
�
�n�W��p�j`1pM�1�1�    P�ON_TextExtra    D90490A5-DB86-49f8-BDA1-9080B1F4E976    ON_DimensionExtra   8AD5B9FC-0D5C-47fb-ADFD-74C28B6F661E    ON_Annotation2  8D820224-BC6C-46b4-9066-BF39CC13AEFB    ON_LinearDimension2 BD57F33B-A1B2-46e9-9C6E-AF09D30FFDDE    ON_RadialDimension2 B2B683FC-7964-4e96-B1F9-9B356A76B08B    ON_AngularDimension2    841BC40B-A971-4a8e-94E5-BBA26D67348E    ON_TextEntity2  46F75541-F46B-48be-AA7E-B353BBE068A7    ON_Leader2  14922B7A-5B65-4f11-8345-D415A9637129    ON_TextDot  74198302-CDF4-4f95-9609-6D684F22AB37    ON_OrdinateDimension2   C8288D69-5BD8-4f50-9BAF-525A0086B0C3    ON_AngularDimension2Extra   A68B151F-C778-4a6e-BCB4-23DDD1835677    ON_AnnotationTextFormula    699FCC42-62D4-488c-9109-F1B7A37CE926    D�0�0��:0���И�p� ��`������W� �ON_Linetype consecutive segments have length zero.
 ON_Linetype consecutive segments have same type.
   ON_Linetype segment has invalid m_seg_type.
    ON_Linetype segment has negative length.
   ON_Linetype bogus single segment linetype - type != stLine
 ON_Linetype bogus single segment linetype - length <= 0.0 (it must be > 0)
 ON_Linetype m_segments.Count() = 0
 line    space   invalid Pattern = ( Pattern length = %g
    Segment count = %d
 ON_Linetype 26F10A24-7D13-4f05-8FDA-8E364DAF8EA6        ������������������������� ������� �h�Я��<�����2P2 �����@����@��@���������� �`�bool value
 integer value
  number value
   point value
    vector value
   xform value
    rbg(%d,%d,%d)   color value
    uuid value
 string value
   object id:  objref value
   polyedge value
 ��P�p��p���0�p������������    ��� ���������p�����������    h�p�������� ����p���������    �� � ��Р�p�����p��������     ���������������p�������    L� �@�� �� �������p������    ������� �������p����������    ��@�`��0�@� ��������p�����0�����@� �rp�`�0�@��W� �Value ID %d:
   none
   Values:
    Descendant ID:
 No descendants.
    Antededent ID:
 No antededents.
    Record type: %s
    history parameters  feature parameters  Record ID:  Version %d
 Command ID:         |���0��P�`�P��������������    ��@����p������������������    �@�������� ��������������ON_HistoryRecord    ECD0FD2F-2088-49dc-9641-9CF7A28FFA6B    `������ @� ��������W� ������Userdata extension of ON_Hatch (contains basepoint) Loop type is invalid.
  2d loop curve has non-zero z coordinates
   Loop curve is not valid
    2d loop curve is NULL
  2d curve:
  2d curve: null pointer
 Inner hatch loop
   Outer hatch loop
          ���￰�@��2 3��������<�Line[%d] is not valid.
 Line type patetern with no lines.
  Type field not set correctly.
  Loop[%d] is not valid
  Loop[%d] is NULL
   Plane is not valid
 %lf 
Dash count = %d:    offset =    base =     ON_HatchLine: angle = %lf radians ( %lf degrees)    Line count = %d
    Description: %ls
   fill type: Solid    fill type: Lines    fill type: Gradient Hatch pattern -     @�������  ��`�������� � �@���@���
�
�n�W��pq��Loop count = %d
    Plane z axis: %g, %g, %g
   Plane y axis: %g, %g, %g
   Plane x axis: %g, %g, %g
   Plane origin: %g, %g, %g
   Base point: %g, %g, %g
 Pattern scale: %g
  Pattern rotation: %g
   Hatch: Pattern index: %d
   ��@���`  ��`�`� ����W  �ON_HatchExtra   3FF7007C-3D04-463f-84E3-132ACEB91062    ON_HatchPattern 064E7C91-35F6-4734-A446-79FF7CD659E1    ON_Hatch    0559733B-5332-49d1-A936-0532AC76ADE5    ���  � ��`�`��W� �group name = "%ls"
 group index = %d
   ON_Group    721D9F97-3645-44c4-8BE6-B2CF697D25CE          �(��
�	����p�@ 
�
�
��� � @!`!0 @ ���W�@�!� r@��
�
�n���k�p�B! k�!p"�" #�Y@#�#%$p&�#�&p' '�'��'`�( !	�B k )P)p)�)ON_OffsetSurface    00C61749-D430-4ecc-83A8-29130A20CF9C        ���*�+ @!`!0 @ ���W�@�!� r@��
�
�n���k�p�B! k�!p"�" #�Y@#�#%$p&�#�&p' '�'��'`(�( !	�B k )P)p)�)ON_SurfaceProxy uses %x
    4ED7D4E2-E947-11d3-BFE5-0010830122F0        $� ,�MpO �/@0P.`.`0�0�W� � �@P r@ 2�
�
�n���k�p�B��@E�4@Q�r 5�Y�r�5 ^�Z6���06�6�6�6�7p9�;p>�Q`A DkkON_PlaneSurface
    .\opennurbs_planesurface.cpp    ON_PlaneSurface::GetNurbForm    ON_PlaneSurface::GetNurbForm - using invalid surface.       x�@,@U U �/�U�K�K�K`L�J� � �@P r@ 2�
�
�n���k�p�B��@E�4@Q�r 5�Y�r�5 ^�Z6���06�6�6�6�7p9�;p>�Q`A DkkPlane surface
  Plane ID =  View IDs =
 Enabled = %d    Clipping plane surface
 ON_PlaneSurface 4ED7D4DF-E947-11d3-BFE5-0010830122F0    ON_ClippingPlaneSurface DBC5A584-CE3F-4170-98A8-497069CA5C36    ���W�W�l ����;����W� ����� r@�p�
�
�n���k�p�B�� k���X�����Y��@Z ^�Z�a v��@m�y�������a !	�B k�a�Wkk      �>      �?������<�4ED7D4E1-E947-11d3-BFE5-0010830122F0      point   NO point array
   ON_PointGrid size = %d X %d
    0� �@�Ќ ��@�`����� � ���0�@��0/0/ ��W��pqON_PointGrid    4ED7D4E5-E947-11d3-BFE5-0010830122F0    �� ���� ����`�0����� � �`�@�@��0/0/���W��pq (hidden)   , normal =  point[%2d]:     ON_PointCloud: %d points
   ON_PointCloud   2488F347-F8FA-11d3-BFEC-0010830122F0    ON_Annotation has m_type = ON::dtNothing.
  ON_Annotation: ....
    % c < >     < > % c     ��`�P�@� @���`��� ���� � ��8 r@�0/0/��W��pqON_AnnotationTextDot.m_text is empty
   ON_AnnotationTextDot "%ls" at   $���Ф�� �� �`�P��� �� � �� r@p��
�
�n�W��pqON_AnnotationArrow has m_head=m_tail.
  ON_AnnotationArrow:     �u �<�7�t���W@�  �P�`�p� � �� � �p� r@��
�
�n�W��pq��`�P�    ��P.5�_��P��`�  �P�`�p� � �� � �p� r@��
�
�n�W��pq��`�0�    ���0���  �P�`�p� � �� � �p� r@��
�
�n�W��pq��`�P�    l�Ж����  �P�`�� � �� � �p� r@��
�
�n�W��pq��`�@�    ��� ��  �P�`�К� �� � �p� r@��
�
�n�W��pq��`�P�    �P�`��  �P�`�p� � �� � �p� r@��
�
�n�W��pq��`�P�ON_Annotation   ABAF5873-4145-11d4-800F-0010830122F0    ON_LinearDimension  5DE6B20D-486B-11d4-8014-0010830122F0    ON_RadialDimension  5DE6B20E-486B-11d4-8014-0010830122F0    ON_AngularDimension 5DE6B20F-486B-11d4-8014-0010830122F0    ON_TextEntity   5DE6B210-486B-11d4-8014-0010830122F0    ON_Leader   5DE6B211-486B-11d4-8014-0010830122F0    ON_AnnotationTextDot    8BD94E19-59E1-11d4-8018-0010830122F0    ON_AnnotationArrow  8BD94E1A-59E1-11d4-8018-0010830122F0    h�p�����  �����0���0����p1��`�@@�0/0/�n�W��pq.\opennurbs_nurbsvolume.cpp m_varient = %d - should be 1, 2, or 3
  Control object:
    Varient: %d
    ����p����
  CV[%2d][%2d]      ON_NurbsCage dim = %d is_rat = %d
        order = (%d, %d, %d) 
            cv_count = (%d, %d, %d) 
   ON_NurbsCage::Create - invalid orders   ON_NurbsCage::Create - invalid cv counts    ON_NurbsCage::Create - invalid is_rat   ON_NurbsCage::Create    ON_NurbsCage::Create - invalid dim  ON_NurbsCage::GetBBox   ON_NurbsCage::GetBBox - invalid input   ON_NurbsCage::Read - invalid dim    ON_NurbsCage::Read - invalid order0 ON_NurbsCage::Read - invalid order1 ON_NurbsCage::Read - invalid order2 ON_NurbsCage::Read - invalid cv_count0  ON_NurbsCage::Read - invalid cv_count1  ON_NurbsCage::Read - invalid cv_count2  ON_NurbsCage::Read - invalid is_rat ON_NurbsCage::Read  ON_NurbsCage::Read - old code unable to read new version of chunk        �����P���������@�p�p�������P�@���
�
�n�0��pqON_NurbsCage    06936AFB-3D3C-41ac-BF70-C9319FA480A1    ON_MorphControl D379E6D8-7C31-4407-A913-E3B7040D034A    P�0� �p� �@�P������p���� �������@���
�
�n�W��pqON_DetailView   C8C66EFA-B3CB-4e00-9440-2AD66203379E    ������p� ������������p�� �P�`���@��0/0/���W��p0p��p��� !	������=���= � ��]
�>�p��W�W`IPh���P�P�p�p����� D ^
 ^
length = %g
    
end =  start =     ON_LineCurve:  domain = [%g,%g]
    ON_LineCurve::Split - input right_side not an ON_LineCurve* .\opennurbs_linecurve.cpp   ON_LineCurve::Split ON_LineCurve::Split - input left_side not an ON_LineCurve*  ON_LineCurve    4ED7D4DB-E947-11d3-BFE5-0010830122F0        �����p ��������p��@�!�P]@��
�
�n�W��p0p 0 !	�<�=�. ��%p�>p���P��A�AP�@G� ���ON_CurveProxy.m_this_domain is not increasing.
     ON_CurveProxy.m_real_curve_domain is not included m_real_curve->Domain().
  ON_CurveProxy.m_real_curve_domain is not increasing.
   ON_CurveProxy uses %x on [%g,%g]
   4ED7D4D9-E947-11d3-BFE5-0010830122F0    ��(�0�1 p*0+�(�P+�+p�� � - -P]@@-�
�
�-�W��p0p���-�]
 !	�<@.`.=�.�.�. !	0/�>�/�a�/�/`IPh�/�A�A�1�@G�]
@0�WHH    ON_CurveOnSurface::IsValid() m_c3 and m_s have different dimensions.    .\opennurbs_curveonsurface.cpp  ON_CurveOnSurface::IsValid  ON_CurveOnSurface::IsValid() m_c2 is not 2d.    ON_CurveOnSurface 
 ON_CurveOnSurface::GetNurbForm  TODO - finish ON_CurveOnSurface::GetNurbForm(). ON_CurveOnSurface   4ED7D4D8-E947-11d3-BFE5-0010830122F0        \��8�K�L @=�=; ;�>0?p�� �0��; �@=�
�
�n�W��p0p��p@�?�L0@���@=��= !	 !	�@�>@A�A�A�A`IpN�ApMP�A0E�F�R�h�I�i�jON_ArcCurve m_arc is not valid
     ON_ArcCurve - m_t=(%g,%g) - it should be an increasing interval.
   
radius = %g
   center =    ON_ArcCurve:  domain = [%g,%g]
       `@���8�K�L @=�=; ;�>�Ip�� �0��; �@=�
�
�n�W��p0p��p@�?�L0@���@=��= !	 !	�@�>@A�A�A�A`IpN�ApMP�A0E�F�R�h�I�i�j          �?      �?      �?�(���!@      �<tbez>=-ON_ZERO_TOLERANCE && tbez<=1+ON_ZERO_TOLERANCE is false       �?.\opennurbs_arccurve.cpp    ON_Arc::GetNurbFormParameterFromRadian  descrim>=0 is false ON_ArcCurve CF33BE2A-09B4-11d4-BFFB-0010830122F0    ON__OBSOLETE__CircleCurve   CF33BE29-09B4-11d4-BFFB-0010830122F0    ��l�WPq ���`����W� ����� r@�p�
�
�n�W��pq4ED7D4DA-E947-11d3-BFE5-0010830122F0    �������?I   ��s�{w  t0w`�@t�y�W� �font linefeed ratio = "%g"
 font is underlined = "%d"
  font is italic = "%d"
  font weight = "%d"
 font face name = "%ls"
 font name = "%ls"
  font index = %d
    A r i a l   .\opennurbs_font.cpp    ON_Font::Read   ON_Font::Read - get newer version of opennurbs  ON_Font 4F0F51FB-35D0-4865-9998-6D2C6A99721D    Userdata extension of ON_DimStyle   h�0�@��� ���`�p�P��W  ���]     [     dimstyle name = "%ls"
  dimstyle index = %d
    ��`|�� � @� ��}��}@�W� ������ON_DimStyleExtra    513FDE53-7284-4065-8601-06CEA8B28D6F    ON_DimStyle 81BD83D5-7120-41c4-9A57-C449336FF12C        �@��WП ��P�`����W  ���������������size of image = %d bytes
   bits per pixel = %d
    height = %d pixels
 width = %d pixels
  P������ p�P�`�p� ��W  �0�@���P�������ON_WindowsBitmap is not valid
      ��P��`� p�P�`������W  �0�@���P�������.\opennurbs_bitmap.cpp      ON_WindowsBitmap::ReadCompressed() image bits buffer size mismatch
 ON_WindowsBitmap::ReadCompressed    ON_WindowsBitmap::ReadCompressed() buffer size mismatch
        �������� ��P�`��`��W  ��W�W�W�W�W��ON_EmbeddedBitmap m_buffer = 0
 ON_Bitmap   390465E9-3721-11d4-800B-0010830122F0    ON_WindowsBitmap    390465EB-3721-11d4-800B-0010830122F0    ON_EmbeddedBitmap   772E6FC1-B17B-4fc4-8F54-5FDA511D76D2    ON_WindowsBitmapEx  203AFC17-BCC9-44fb-A07B-7F5C31BD5ED9    D  ���<�� �      .@      4@      <@      L@     �Q@     �F@      ^@     @j@     �o@     �P@     �k@     �~@     ��@     ��@     �V@     �v@     H�@     H�@     v�@     Ъ@      ^@     ��@     p�@     �@     H�@     X�@     #�@      c@     ��@     �@     ��@     !�@     �@    �]�@    ���@     �g@     Б@     �@     H�@     ��@     ��@     ��@    ��A    ��A     �l@     �@     ��@    ���@    P7�@    ��A    h�A    0\A    �#A    0�%A     @q@     ��@     ��@     ��@     n A    �A    �q&A    p�3A    (�=A    HCA    ��DA     Pt@     P�@     3�@    @�@    �A    $A    ��7A    ��GA   �=CTA    y]A   ��kbA    k�cA     �w@     ��@    ���@    ���@    ��A    (2A   ���GA    YZA   ��iA   @�ztA   �/}A   ��ځA   �!�A     0{@     ��@    @��@    PeA    �"A    X?A   @�SVA   ��IkA   p5�|A    _�A   � ��A   ����A   ��U�A   ��}�A      @     `�@     ��@     �A    ��+A    �IA   ��dA    ڿzA   �ÎA   �ÞA   ���A    ���A   P��A   0��A   #���A     ��@     `�@     ��@    ��A    ��4A    ��TA   ��PqA   ���A   0mC�A   `��A   ��W�A   H���A   6���A   H���A  �
�k�A  �) c�A     ��@     �@     ��@    �A    ��=A    �_A   @��|A   �r�A   �*M�A   ����A   �Ŧ�A   <{7�A   ��H�A   6���A  �vT9�A  �� B   �\� B     ��@     z�@    p�@    آA   ��EA    <hA    �Q�A   p�n�A   <X-�A   lO��A  �Y,�A  �Y,�A  �}�B   �H�B  xPl�B  P���B  ���EB  p�{u B     `�@     L�@    �O�@    �$A    �HMA   ���qA   ��U�A   �XL�A   �"C�A   Li9�A  ��	��A   G�iB  ����B  @<�"B  $�D-B  ��ܨ4B  ��e:B  Г
�>B  ��%@B     �@     l�@    �S�@    ��)A   ��TA   ���yA   ��#�A   �ē�A  @��A   ܅��A  ���B  @�#�B  �+n�(B  `�U�6B  \`bCB  zP��MB ��p�TB  t�xZB  �p�]B  �תT_B     ��@     ��@    8� A    8�0A    ��ZA   ��E�A   � �A   � �A  @)�|�A  �?��A  �i�B  @"�,(B  o��:B  o��JB ��ԈAXB  k���cB �����mB �fN�tB `��a�yB  ͑�I}B �$a�~B     ,�@     ��@    ��A    ��4A   `��aA   @ƅ�A   �	�A  �ڶj�A  �z_�A  ��a�B  nЁ"B  s��7B �"l��KB  Xs��]B @�o4�lB �j5vyB p�����B �r-�9�B ���g�B ����B�B x�{��B �����B     ��@     ��@    ��A    � :A    �ggA   @���A   ��}�A   t���A  �w�]�A  ��B  �x�80B  躵uFB  �)#\B  l�oB x���g�B  ����B @��З�B @�|���B Pu(q�B �NpK�B p�_8�B ���'�B _�:T�B     $�@     $�@    �A    4*@A   �!OnA   �uЗA    �A  �L���A  �44"B  `��d!B  ��C<B  2sէTB �]�~KkB ��-`�B \���B \���B ?-jk�B �Tto��B �'��n�B h�@��B V�M�-�B �.���B �-��B ^����B     ��@     ��@    �A    �CA   �WjsA   ���A   im�A   �Gi�A  �L�wB  ��� ,B  �HB  �>8{bB ����yB �Y��M�B ���٢B ,�����B y��g�B ��V�\�B�݂Bڥ�B l�{���B ^�Œ��B γj��B@�Cַ<�B g�H%�B���0�B.\opennurbs_math.cpp    ON_GetPolylineLength    ON_GetPolylineLength: Zero weight   .\opennurbs_knot.cpp    ON_KnotVectorSpanCount  NULL knot[] passed to ON_KnotVectorSpanCount.   ON_GetKnotVectorSpanVector  NULL knot[] or s[] passed to ON_KnotVectorSpanCount.    ON_IsKnotVectorPeriodic ON_IsKnotVectorPeriodic(): illegal input    ON_SetKnotVectorDomain - invalid input  ON_SetKnotVectorDomain  ON_SetKnotVectorDomain - invalid input knot vector  Knot vector order = %d but knot[%d]=%g >= knot[%d]=%g
  Knot vector must be increasing but knot[%d]=%g > knot[%d]=%g
   Knot vector cv_count=%d and knot[%d]=%g >= knot[%d]=%g (should have knot[cv_count-2] < knot[cv_count-1]).
  Knot vector knot[%d]=%g is not valid.
      Knot vector order=%d and knot[%d]=%g >= knot[%d]=%g (should have knot[order-2] < knot[order-1]).
   Knot vector knot array = NULL.
 Knot vector cv_count = %d (should be >= order=%d )
 Knot vector order = %d (should be >= 2 )
   ON_MakePeriodicKnotVector(): illegal input  ON_MakePeriodicKnotVector(): illegal input degree=1, cv_count<4 ON_MakePeriodicKnotVector(): illegal input degree=2, cv_count<5 ON_MakeKnotVectorPeriodic       ON_MakePeriodicKnotVector(): illegal input degree>=3, cv_count<2*degree ON_InsertSingleKnot() - illegal knot input  ON_InsertSingleKnot ON_InsertSingleKnot() - illegal cv input    ON_InsertKnot(): out of memory  ON_InsertKnot(): requested knot_value at end of NURBS domain    ON_InsertKnot(): requested knot_value at start of NURBS domain  ON_InsertKnot(): requested knot_multiplicity > degree   ON_InsertKnot   ON_InsertKnot(): illegal input  .\opennurbs_evaluate_nurbs.cpp  ON_EvaluateNurbsDeBoor  ON_EvaluateNurbsDeBoor(): knots[degree-1] == knots[degree]  �Z�!@.\opennurbs_zlib.cpp    ON_BinaryArchive::WriteDeflate  ON_BinaryArchive::WriteDeflate - z_deflate failure  ON_BinaryArchive::ReadInflate   ON_BinaryArchive::ReadInflate - z_inflate failure   1.2.3   ON_BinaryArchive::ReadCompressedBuffer  ON_BinaryArchive::ReadCompressedBuffer() crc error  .\opennurbs_objref.cpp  ON_ObjRef::DecrementProxyReferenceCount ON_ObjRef::DecrementReferenceCount() *m__proxy_ref_count <= 0   � �{ {�{�{`���p� �r�0��p�0��W� ������M e s h   N - g o n   l i s t   ON_MeshNgonUserData 31F55AA3-71FB-49f5-A975-757584D937FF    ON_Brep::NewLoop unable to make 3d edge curve.  Bad edge information passed to ON_Brep::NewFace.    Bad vertex index passed to ON_Brep::NewFace.    Bad edge index passed to ON_BrepNewFace.    ON_Brep::NewFace(ON_Surface*,...) error: Bad edge vertex informtion.    .\opennurbs_brep_tools.cpp  ON_Brep::NewOuterLoop       ON_Brep::NewFace(ON_Surface*,...) error: Edge and vertex informtion do not match.   ON_Brep::ReadOld201() - trouble reading render/analysis meshes  ON_Brep::ReadOld200 - trim.m_trim_index out of range.   ON_Brep::ReadOld201 - trim.m_ei out of range.   .\opennurbs_brep_io.cpp ON_Brep::ReadOld200 ON_Brep::ReadOld200 - trim.m_trim_index out of synch.   ON_BrepTrimArray::Read  Invalid value of m_trim_index   B r e p   R e g i o n   T o p o l o g y     lP����� �r�`��� ��W� ��@�P����� @���0�p�H�� ��� �r�`�0����W� ������0�`������0�`�0`���0�`�|`���0�`�    � ����� @�������0��W� �0���p�ON_BrepRegionTopologyUserData   7FE23D63-E536-43f1-98E2-C807A2625AFF    ON_BrepFaceSide 30930370-0D5B-4ee4-8083-BD635C7398A4    ON_BrepRegion   CA7A0092-7EE6-4f99-B9D2-E1D6AA798AA1        Attempt to seek to a position that is too large for 64-bit unsigned int storage.    Attempt to seek before start of buffer. .\opennurbs_embedded_file.cpp   ON_Buffer::Seek Invalid origin parameter    ON_Buffer::Copy Attempt to copy corrupt source. corrupt buffer - list of segments is too long.  corrupt buffer - segments contain more bytes than m_buffer_size.    corrupt buffer - empty segment buffer.      corrupt buffer - previous segment's position1 !- segment's position0.   corrupt buffer - first segment has non-zero value for position0.    ON_Buffer::CRC32    corrupt buffer - segment's position values are invalid. ON_Buffer::SetCurrentSegment    Corrupt ON_Buffer   ON_Buffer::Write    size parameter > 0 and buffer parameter is null.    Uncompressed buffer - m_file_size != m_buffer.Size(0)   m_buffer_crc != m_buffer.CRC32(0)   m_buffer is not valid.  ON_Buffer::ChangeSize   Corrupt ON_Buffer.      The buffer contents were corrupted during, writing, storage or reading. ON_Buffer::ReadFromBinaryArchive    corrupt archive  %�% 0�`���"�W� �ON_EmbeddedFile 1247BEC9-D9A9-46B3-900F-39DE7A355BD3    h�	�� �  �  deflate 1.2.3 Copyright 1995-2005 Jean-loup Gailly             `6    @8    @8      @8    �;      �;  � � �;   �  �;  �  �;   �;1.2.3   `   P   s   p  0  	� 
  `     	�     �  @  	�   X    	� ;  x  8  	�   h  (  	�    �  H  	�   T   � +  t  4  	�   d  $  	�    �  D  	�   \    	� S  |  <  	�   l  ,  	�    �  L  	�   R   � #  r  2  	�   b  "  	�    �  B  	�   Z    	� C  z  :  	�   j  *  	�  
  �  J  	�   V   @  3  v  6  	�   f  &  	�    �  F  	� 	  ^    	� c  ~  >  	�   n  .  	�    �  N  	� `   Q   �   q  1  	� 
  a  !  	�    �  A  	�   Y    	� ;  y  9  	�   i  )  	�  	  �  I  	�   U   +  u  5  	�   e  %  	�    �  E  	�   ]    	� S  }  =  	�   m  -  	�    �  M  	�   S   � #  s  3  	�   c  #  	�    �  C  	�   [    	� C  {  ;  	�   k  +  	�    �  K  	�   W   @  3  w  7  	�   g  '  	�    �  G  	� 	  _    	� c    ?  	�   o  /  	�    �  O  	� `   P   s   p  0  	� 
  `     	�     �  @  	�   X    	� ;  x  8  	�   h  (  	�    �  H  	�   T   � +  t  4  	�   d  $  	�    �  D  	�   \    	� S  |  <  	�   l  ,  	�    �  L  	�   R   � #  r  2  	�   b  "  	�    �  B  	�   Z    	� C  z  :  	�   j  *  	�  
  �  J  	�   V   @  3  v  6  	�   f  &  	�    �  F  	� 	  ^    	� c  ~  >  	�   n  .  	�    �  N  	� `   Q   �   q  1  	� 
  a  !  	�    �  A  	�   Y    	� ;  y  9  	�   i  )  	�  	  �  I  	�   U   +  u  5  	�   e  %  	�    �  E  	�   ]    	� S  }  =  	�   m  -  	�    �  M  	�   S   � #  s  3  	�   c  #  	�    �  C  	�   [    	� C  {  ;  	�   k  +  	�    �  K  	�   W   @  3  w  7  	�   g  '  	�    �  G  	� 	  _    	� c    ?  	�   o  /  	�    �  O  	�    A @ !  	 � @   �  a ` 1 0 � @         	  
             incorrect length check  incorrect data check    invalid distance too far back   invalid distance code   invalid literal/length code invalid distances set   invalid bit length repeat   invalid literal/lengths set too many length or distance symbols invalid code lengths set    invalid stored block lengths    invalid block type  header crc mismatch unknown header flags set    incorrect header check  invalid window size unknown compression method                                                                                                   	
                                                                 	   	   
   
                                                                                                    �  L  �  ,  �  l  �    �  \  �  <  �  |  �    �  B  �  "  �  b  �    �  R  �  2  �  r  �  
  �  J  �  *  �  j  �    �  Z  �  :  �  z  �    �  F  �  &  �  f  �    �  V  �  6  �  v  �    �  N  �  .  �  n  �    �  ^  �  >  �  ~  �    �  A  �  !  �  a  �    �  Q  �  1  �  q  �  	  �  I  �  )  �  i  �    �  Y  �  9  �  y  �    �  E  �  %  �  e  �    �  U  �  5  �  u  �    �  M  �  -  �  m  �    �  ]  �  =  �  }  �   	 	 � 	 �	 S 	 S	 � 	 �	 3 	 3	 � 	 �	 s 	 s	 � 	 �	  	 	 � 	 �	 K 	 K	 � 	 �	 + 	 +	 � 	 �	 k 	 k	 � 	 �	  	 	 � 	 �	 [ 	 [	 � 	 �	 ; 	 ;	 � 	 �	 { 	 {	 � 	 �	  	 	 � 	 �	 G 	 G	 � 	 �	 ' 	 '	 � 	 �	 g 	 g	 � 	 �	  	 	 � 	 �	 W 	 W	 � 	 �	 7 	 7	 � 	 �	 w 	 w	 � 	 �	  	 	 � 	 �	 O 	 O	 � 	 �	 / 	 /	 � 	 �	 o 	 o	 � 	 �	  	 	 � 	 �	 _ 	 _	 � 	 �	 ? 	 ?	 � 	 �	  	 	 � 	 �	    @     `    P  0  p    H  (  h    X  8  x    D  $  d    T  4  t    �  C  �  #  �  c  �                       
                	                         								















   		

                            
                         (   0   8   @   P   `   p   �   �   �   �                                              0   @   `   �   �      �                               0   @   `      �0w,a�Q	��m��jp5�c飕d�2�����y�����җ+L�	�|�~-����d�� �jHq���A��}�����mQ���ǅӃV�l��kdz�b���e�O\�lcc=���� n;^iL�A`�rqg���<G�K���k�
����5l��B�ɻ�@����l�2u\�E���Y=ѫ�0�&: �Q�Q��aп���!#ĳV���������(�_���$���|o/LhX�a�=-f��A�vq�� Ҙ*��q���俟3Ը��x4� ��	���j-=m�ld�\c��Qkkbal�0e�N b��l{����W���ٰeP�긾�|�����bI-��|ӌeL��Xa�M�Q�:t ���0��A��Jו�=m�Ѥ����j�iC��n4F�g�и`�s-D�3_L
��|�<qP�A'�� �%�hW��o 	�f���a���^���)"�а����=�Y��.;\���l�� �������ұt9G��wҝ&���sc�;d�>jm�Zjz���	�'� 
��}D��ң�h���i]Wb��ge�q6l�knv���+ӉZz��J�go߹��ﾎC��Վ�`���~�ѡ���8R��O�g��gW����?K6�H�+�L
��J6`zA��`�U�g��n1y�iF��a��f���o%6�hR�w�G��"/&U�;��(���Z�+j�\����1�е���,��[��d�&�c윣ju
�m�	�?6�grW �J��z��+�{8���Ғ�����|!����ӆB������hn�����[&���w�owG��Z�pj��;f\��e�i�b���kaE�lx�
����T�N³9a&g��`�MGiI�wn>JjѮ�Z��f�@�;�7S���Ş��ϲG���0򽽊º�0��S���$6к���)W�T�g�#.zf��Ja�h]�+o*7������Z��-    A1�b62�S-+�ldE�w}��ZVǖAO���I��ъ�������O��M~���-�����Q�J#�S�p�x�A�aU׮.�7׵����Y��� ���-���6�]]w�ll��?AԞZ͢$����� F��aw����������$���e��ڪ�]]�FD(�koi�pv�k19�Z* ,	m8�6F߲]�qTp�0ek���*���1�u��4��������yީ%8�<�y�s�H�j}�A<*�XOy�D~b�-O��T���@����#���8�Š8L��!���
Ζ�	 �\H1�E�b�n�S�wT]��l���?�����P�������������\�br�yk޵T@��OYX#�p8$�A#=�k�e�Z�|%	�Wd8�N���⟊!̧3`��*��$���?�-��l�	��$H��S�)F~�hwe��y?/�H$6t	5*�SK��HRp�ey1�~`�������|���=����6�����xT��9e��K��;
��"���	�ˮO]�_l�F�?�m��tCZ�#A��pl��Aw�G�6��-�ŵ �����Aq[�Zh��wC��lZO-_~6�-'� > ��S1���b���S�����W��Ĕ���Ֆ�������k�1�*�*��ykʬHp�o]�.*F��6�f��cT�T"e�M���©g��0&��)��������:���{��ϼk���Z��>	��8���$,�52F*sw1��pH��kQ6�Fzw�]cN������̵������J��#���p���A��F]#l8�?1�(B�Og�T~��yU��bL�8�^�#����ܖ� T�Z1O��bb��Sy�O�IV~�P�-�{��b��-R��4���٠��~^��eGn�Hl/�Su�6:�	#jT$+e?�y���H��f��'*�������b���#��ٽ��Ч?��&~��?�$�p��i;F�Bzw�[�ke��Z~�7	S�v8H���	���3�?�r�$�    7j�nԄY�Fܨ	����|��O�Q�;�օ���Ud�	S��
-�
=G\p�&G��w�)`�/�a��߫��i��5����&��LsZ<#0�z��M�z�FM8�,�9���;��:<�D?��>R:�<eP=X^6o}�76��5�4��W1�Օ0�k�2�3��k$���%�1�'�[-&LMb#{'�""�� �$!(�x*޺+F`�)q
>(�q-�v�,���.��7/���p��Xq�Ys�3�r%�w+OQvr�tE��ux܉~O�K}!b�|�t�y�Bxʠz���{�.�l�D~m��8o��nl��k[�wjR1h58�i�b?mcf�+aQ��`�צe�dd�"f�i�g ��H�INSKyu�J�c�O�	N��ZL�ݘM���F��G�N@E�$�DD2�AsX@*�IB��CPh�Tg3U>�uW	ַV���S��:R�|P�~�Q�9�Z�S [��fY���X4��]�)\ZEo^m/�_�5�q���ϱ�٥s�\�<�k���2g��z�8J&� ��V���a�`���/�ӈ��6��\i��������l���U�,�z��BĞ�u�\�H� ����&=��WF�A	��+��������O�`]x�W7�����9�>ۼ�qދ����!���K7��k��f�ֶ��ԁ�-��b�3Π�jp��]$��^�'���~*��I@��VW��<�â��������M˟ŏ��{����tD�Cm�����-��@���w�m�.B+�(铜>���Td���"�ŀ���Ǽ�ϭ~��8��y��$o��w�J�1�}��05��_K�^��i�Ϗ은���B��I��#ƈ�d���X�����܁T̓�c�Q�:�rՆ��⩗� ��f��n��|x�K)��o�%ƭ���/�3�vUu�A?���)���C:���|������sĵ����@��͂��Ͳ;��bI�Ue��h"׻_H��S�1�����޼����^Z��4��    eg����	�W�b�2��7�_k%�8ם�(�ŊO}d�o�׸��J��j�3w��VcX�WP�0����q��B��{߭��gCru&o��p��-���?���'��B�s�� ư�Gz>�2�[Ȏ�g;
� ��i8P/_���Y����=ч�e��:�ZO��?(3w����wXR��@h�Q���+�ğ�H*0"ZOW���oI���}�@���mNП5+�#�����*'G��| A�����H�=X�X?�#��1����j�v�ʬ���`��p�^��Y���<�L������~i/�{kHwâ��h�s)�aL�����oD����~Pf�7�VM'�(@��ﰤ���ہ�g9�x�+�n��&;f����?/��X�)T`D�1�ߨM����ߒ���.Fg�Tp'�H�q�/L�0���U�Ec��?k�ǃ�h6�r�y�7]�P�\@�TN%���s����7�@��'>�$�!AxU�����ʰ\3;�Y�^��U�~PG���l!;b	F����2Ȃ��pԞ�(��Q�_V�:1X:�	���n3��m�:���@����/)IJN���v"2���x�+�ٗ K��x.�H���ҥfAj^��y9*O���]��#�kM`~����b���_R�	�7�z�F h�!���1߈�Vc0a��"�j�������6n��S	�Nr�)Υ�{�t��������*F8#v��uf��z`���r��s�"�WG��9���^E�Mvc��΍&D��A�dQy/�4�Aڱ&S�֚�������Eb�iL��Q�<�6'�5���P�..��T&���q]�w�4�.6��I�E�? ���v����\[�Y�I�>U�!�lDa>Ԫ΋�ϩ7~8A�]&�n��v|����o�Y
�����y�K�i��w�\�¹9�~�����$6�6nQ��f��q�>,�o,I�Ӕ��	�渱{I�.�H>�C-Yn����馑gQ���z�t�a�f��    w0��a,�	Q�m�pj��c�5�d��ۈ2yܸ������و	�L+~�|��-����dj� ��qH��A���}m����ԵQ�Ӆ�l�Vdk���b�z�e��\Ocl��=c��;n �Li^�`A�gqr<��K�G����
�k5���B��lۻ�֬��@2�l�E�\u��ϫ�=Y&�0�Q� :��Q���a!���V��#Ϻ�����(��_��ٲ��$/o|�XhL�a��f-=v�A��q�� ���*q����������3xɢ �4�	����j�m=-�dl��c\kkQ�lab�e0��b Nl���{�����We�����P�������|b���-I��|���LeM�aX:�QΣ� tԻ0�JߥA=ؕפ��m����Ci�j4n���g�F�`��D-s3�
L_�|�Pq<'A��� �Wh�% o���f�	�a�^��)�ɘ�И"�ר�Y�=.����\;��l�� ������t�Қ��G9��w��&s���c�d;�mj>zjZ����	��
 �'}����D����hi���bW]�eg�l6qnk���v��+��zZg�J����o������C`����֣�ѓ~8���O��Rѻg�Wg?��H�6K�+گ
L6J�Az`�`�èg�U1n��Fi�y�a���f�%oҠRh�6�w��G"�U&/ź;���(+�Z�\�j�������1,ٞ�[ޮ�d°�c�&uj��m�
�	��6?rg� W��J��z{�+��8�Ҏ��վ|����!�������Bhݳ�ڃn�����&[o�w��Gw�Z��jpf;�\�e���b�iak��l�E�
�x���N�T9�§g&a�`�IiGM>nwۮ�jJ��Z�@�f7�;𩼮S޻��G��0��齽�ʺS��0$�����6���T�W)#�g��fz.�aJ�]h*o+���7���Z�-�    1A26b�+-S�dl�}w�EVZ��OA���ي�»I������ˬ�O��~M��-����J�QS�#x�p�a�A�.��U7����������Y� ��-�۩6˚�w]]�ll�A?��Z���$���㧲F ��wa��������ރ$�Ųe]]��DF��ok�(vp�i91k� *Z�	,8m�F6��]��pTq�ke0�*���1¶��u��4������%��y<��8s�y�j�H�A�}X�*<�yO�b~D�O-��TƔ���@�#胿8��8��!��L
������\� 	E�1Hn�b�w�Sʺ�]T��l��?֑���טP�̩������˓rb�\ky�@T��YO��X#$8p�=#A�e�k�|�Z�W�	%N�8d������3��!*��`�$᯴?���-�	�l�H$��S��~F)�ewh/?y�6$H�	t*5KS��RH��ye�p`~�1������¿�Б|�ˠ=��6������Tx��e9;��K"��
	����ˈ_�]OF�lm�?�t���ZC�A#�lp��wA��6�G�-�� �ż��qA�hZ�[Cw�Zl��-O6~_'-�> ݹ� ��1S��b���S�������W�§��ٖծ�����1�k�*�*�ky��pH��]o�F*.f�6���T�TcM�e"����¤0��g)��&�Ů��ޟ����:���{��k���Z���	>��8,$�5�*F21wsHp�Qk��zF�6c]�w���N����̵��ׄ���J��#��pȄ�A�#]F8l1?�(�gO�B~T�Uy��Lbˁ�8��#�^�������T �O1Z�bb��yS�I�OP�~V{�-�b��-��4��R�����^~��Ge­lH�nuS�/:6�#	�$Tj?e+��y䏼H���f��*'�˼��Ѝ����b���#�����&��??��~p�$�i��B�F;[�wz�ek��~Z��S	7�H8v�	������?�3�$�r    �j7��nF�Y	������|�O�Q��;����U��	�dؓS
�-
\G=&�p��G�w`)/��a����i��5������&�sL�<Z�0#��zz�M8MF�9�,�;ɒ�:��?D�<>��<�:R=Pe6^X7�}o5��64�1W��0�ճ2�k�3�$k�%���'�1�&-[�#bML"�'{ �"!$�*x�(+��)�`F(>
q-q�,�v�.�Ț/7��p���qX��sY�r�3�w�%vQO+t�ru՛E~��xK�O}|�b!y�t�xB�z��{���l�.�m~D�o8��n���k��ljw�[h1Ri�85b�cm?a+�f`��Qe���dd��f"�g�i�H�� I�KSNJ�uyO�c�N	�LZ��M�ݥFĚ�G�E@N�D�$�A�2D@XsBI�*C��T�hPU3gWu�>V��	S���R:��P|�Q�~�Z�9�[ S�Yf�X���]�4\)�^oEZ_�/m�5���q�����s���<�\���k�g2�z�&J8�� 좞V�`�a�/������6��i\����������l��U��,��z���B�\�u� �H���=&�FW�	A���+������O���x]`غ7W����>�9�q��߳����!��7K��k�֩f���ض�-���b�Ѡ�3��pj�$]�^�Ĝ�'��*~�@I�WV�Õ<��ӂ����M��ʏş��{����Dt͆mC�����-���@�m�w�+B.��(��>��dT��"����ş����~�Ϝ8���y���o$�w�1�J���}��50�K_��^�ϋi����B�ۉI���#���d��X������ф��T�Q�c�:��r��Р� ���fΫ�n���x|�)K�o����%���3�/�uUv��?A��)ġ:C�|��������sд�@����͉�����;�Ib��eU��"h�H_�S����1�ފ�����Z^ھ�4�    ��ge�	ȋ���b�W7��2%k_ܝ�8�Ŵ(�}O�o��d��Jֿ��j����w3XcVPW��0���B��q�{��gǧ�urC��o&��p-?����О��'�s�B�� �zGɠ2�>��[
;g��� �/P8i��_�Y��=嗇e����:�ϏOZw3(?���RXw�@���Q�h�+��H���Z"0*�WOIo�����@�}m��5��N�#�+���'*���GA |􏒨H���X=#�?X1������v�j�ʨ���`�^�p������YL�<���i~��{�/�wHk��s�h�a�)ٸ�LDo�������fP~V�7�'M�@(�������۰9g�+�x��n�;&����f�/?�)�X�D`T�1M�ߦ�Ϻ����F.��T�g�'pq�H��L/����0cE�Uk?��Ӄ���6hy�r�]7�\�P�NT�@��%���s7��@��>'�!�$�UxA��ׯ3\���Y�;U��^GP~����b;!lڇF	�2��p���(�ԐQ����V_:X1:��	�3n����:�m�@����I)/��NJ2"v���+�x ��x��K�H�.���jAf���^O*9y]����#��Mk��~`�bю_޶��	�Rz��7h F�м!���1�0cV�"��a�j������ح�n6	SrN���)��{���t���*���8F��v#��fu`zrϮ��sɛW��"��G��9�E^�vM���c�D&�d�A��/yQA�4S&���ֿ����E���b�Li<�Q��'6ۖ��5..�P&T�������]q4�w�6.��I�?�E��� ���v[\�I�Y��U>�l�!�>aDƋΪ~7���A8n�&]|v������Y�oᡱ
��K�y��i׫w��¡\~�9����$��6�6�Qn�f�>�q�,o�,�ӹI	��散I{�.C�>H�nY-����Qg��̰�t�zf�a���incompatible version    buffer error    insufficient memory data error  stream error    file error  stream end  need dictionary ��t�k4h�X�L�8�(��k4 inflate 1.2.3 Copyright 1995-2005 Mark Adler         	 
         # + 3 ; C S c s � � � �                                    � �         	    ! 1 A a � � � 0@`                                  @ @ string too long invalid string position ��� �֌Unknown exception   _�j8j8csm�               �                          �?      �?3      3            �      0C       �       ��              ������ ������ 3      3             �       �                      �?      �?3      3                      �                     �CorExitProcess  mscoree.dll ..  .   *?  �#�֌bad exception   .mixcrt EncodePointer   KERNEL32.DLL    DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    �`�e+000          �~PA   ���GAIsProcessorFeaturePresent   KERNEL32          �?5�h!���>@�������             ��      �@      �        runtime error   
  TLOSS error
   SING error
    DOMAIN error
  R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:                      �?    ���?     ��?    �D�?    ��?     ��?    @��?    @W�?     �?    ���?    ���?    �w�?    �A�?    ��?    @��?    ���?    �q�?    �?�?     �?    @��?     ��?    �}�?    �N�?    @ �?    ���?    ���?     ��?     m�?    �A�?    ��?    ���?    ���?    ���?     q�?    �H�?     !�?    ���?     ��?    ���?     ��?    �a�?    �<�?     �?     ��?    @��?    @��?    @��?    �g�?    �E�?    @$�?     �?     ��?    ���?    @��?    ���?     b�?    �B�?     $�?    ��?    @��?    ���?     ��?    ���?     r�?    @U�?     9�?     �?    @�?     ��?    ���?    ���?    @��?     {�?    �`�?     G�?    �-�?     �?     ��?    @��?    ���?    @��?     ��?    @��?    �i�?     R�?     ;�?     $�?     �?    ���?    @��?     ��?     ��?    @��?    ���?    @s�?    @^�?    @I�?    @4�?    ��?    @�?     ��?     ��?     ��?    @��?    ���?    @��?     ��?     n�?     [�?    @H�?    �5�?    @#�?     �?     ��?     ��?    @��?    ���?     ��?    ���?    @��?    @��?    @s�?    @b�?    �Q�?     A�?    �0�?    @ �?     �?      �?                          �a���?���F��<=  z1%�?�Vd?E=  ��b�?�6��\�M=  ���?p�9t^�<= �\c�N�?	�ʽ��J= �3���?�/��N=  �b�?DZ.�0=  �Ohe�?�?���0=  ]3��?��`$= @�׹ƻ?X&eB�E= ���rr�?\�3#�.J= ��׌�?��C5= �3:���?Ltm��YE= @�'z+�?�"e���=  tLVv�?p��$��M= `�dH��?h6_~��(= `x��?��Y�O= ���YL�?wJ�Q�\C= ��jU��?�Vш4= �+0��?e���37.= `�2�?�⋱�K= `���I�?)-��W�0=  -�Ƀ�?���*D= ���D��?7Tf(��G= �6	�x�?Y��8= ��%��?�E�<= ��w��?�~�?= �Ґ�C�?]���u�<= P��W��?>#�4�<  ��Xq�?���B�J= �_D��?m��K��F= ��Ԛ�?��s7�E= @�[-�?K>�d�:= ��g��?Z}�=\uI= �s�~Q�?�g:"(�N= �'��?9�~$O1=  ��q�?�n�1��%= p)k� �?v�ʌ�= `�X:��?�q.W�� = Pi���?g���>�M= ��[��?ֲa
��M= �_�3�?֍,�uXO= `Ɏ/��?���1w<= �>'eH�?`�	J�J= x~��? �&= n�`Y�?��˖��C= 0����?�]��/= # �g�?u�P�= �����?���,l�C= �5��q�?ᕎ�	= @Dӳ��?�-[�@= pt�4z�? �فpnJ= ���l��?�i�.Eg�< �y~�?�?�O�^'= (T�t��?�
�x;�;=  �P��?�R�RF= ��&�?X��ɣN= �J��@�?��~��= Ht=c��?Az�U"= ��nB��?U_l�j7= ��]���?q���BD=  �h<�?z�)�t'= �Z�#z�?��0�L= @5��ڿS�OO�F� ��ڿ���ۓ�D� 0���ٿ��= �n�  �W9!ٿ?�j>� 0�"�ؿ�؍� �I� �Q�n0ؿ�Hn&�E� �:�׿E7D���5� ��7�A׿��%@� @���ֿ* ��Z+A� �S��Tֿ�rJ� �D� @ӑ��տ����NT?� �w3�kտr�1�9�  �]��ԿF�K�m�8� �C!`�Կ1y2�Y�� @��Կ*�(<j�  䃝ӿV�CD� p��,ӿ1���n� ��ҿ2�=l�7� 0���IҿO���	x*�  �l@�ѿ2��>�FE� �O�5iѿ���4�Q!� �?:	�п�C	 ��+� pڌX�п��xO,�C�  �"пA��ri<� �q~�_Ͽ�R� v=� �=	~�ο����o6� @m�P�Ϳ	 ���d+� �>��̿9Ȓ���� �[\�˿8�B��'� ����&˿�i�[J� ��Z�Oʿ�b�n�E� �D�E}ɿ�Ugc@� �H	��ȿUZ�d��L�  "� �ǿ=��Dj!�  ��ǿ��Vm�:A� @��`3ƿ�~%�3�  k��cſ�"�7M�  ����Ŀ��p��>� �)%��ÿ\�����B� ��jx�¿#6HQ;� `t�-¿=]P��H0� �;T�a�����ָE�  &�����a-#��K� �V\���Vb���4M� @������U@�  X�x�����55� @���캿D��=� �iI�^��Gי��'7� ��A�Է�U�����N�  ��<N���>Ҫ1� ���Gƴ��O\�C� @��+B���g:IB� @Z�u�������}M� ����:��(T��!1� ���n���]vQ<)8�  h׾o��$�|�f+� ����x��2S��74�  U".���mœFB*� �6�I���KS�_D�   �5��M�-�C�  z1}B����K� G�  �c��?�Of��F�  �L,��s�X4I+�  xm�	w�$��V�cE�                      �?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    @��?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?    ���?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    �
�?    �
�?    @
�?     
�?    �	�?    �	�?    @	�?     	�?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    ��?    ��?    @�?     �?    � �?    � �?    @ �?      �?                          �|)P!?Ua0�		!=   �+34?�2��Q	=  �`��??7;W��J=  `�7�E?��'a %C=  ��MkK?�*��b<=  0ɘP?*�,�z?=  d|S?�K�T'�K=   �R_V?�b���F=  p^�BY?�����E&=  �9&\?�߇�N9=  p��	_?߭Eb2]A=  ���`?��f#I=  ���hb?O2�H`3=  ����c?e2��a�1=  �ԆLe?2���RM=  ����f?A�3�_:=  @�0h?[��2ieO=  ����i?�1r�K=  ���k?����Σ-=  ���l?���̈[8=  �yQ�m?>�|W8A=  �՛ko?�>qݲN=  ���np?z m{M=  t�)(q?m,�S�D=   E`�q?��}e?=  ԩ��r?�}~:f�E=  P��Ss?����&�A=  ��&t?,&��8=  ��t�t?�eѴN�@=  PS�u?^p?o4�0=  �!9v?�W�?N=  <��v?+�#�GYM=  H�w?qC���@=  ��Pex?0&ے=  X��y?���8 =  <8�y?!({=�H=   ���z?�d,G�B=  ��6K{?ҝ��E	M=  �¾|?w�3�1�!=  ��L�|?��^X-F=  �<�w}?0��!�O=  ��y1~?|"į�Q<=  $�~?��k�f@=  �+��?��b�UC=  ��4/�?*�K_�<*=  <��t�?�̍xI=  2�р?wY�V%A+=  ���.�?x+s7�E=  8#o��?�e��fE=  �|R�?Ks޸�E=  T�8E�?�=��(=  ��!��?��)��G=  ���?#F؇K=  V�[�?��C�<  :︃?k�V���I=  ����?����YH=  ���r�?q��4';=  .~�τ?��=�S7=  �'�,�?7���X�#=  4�ԉ�?C��k��7=  bB��?��EpC=  B��C�?'�2xk==  蠆?̸WU�A=  xm�	w�$��V�cE�  ̑ʭv�K��[��7�  �G�Qv�e$�l�F�  ����u��y�ԏ�H�  �gԙu�|��ǣ%I�  ���=u���?FK�  ����t�S'�q	! �  �Yхt�L8|�H�  dw�)t���v�#L�  l&��s���>��D�  �f�qs�g~��7�(�  �7�s���6�uE�  (���r�uv.�E,�  t��]r��L��v�O�  ��r��Ț�p�  �&��q�C �"5�F�  ��zIq�o����O�  �j�p�����O�  |�W�p�Ȯ�/N�  �#D5p�O���/3N�  �^�o��I��!�  `1�n��D�CE�  "Bn��u
^!E�  �WΉm����--�0�  ����l��N���pC�  P&`l����J�  �$ak�����N��  8x�j��[-=�  8R��i�y��~� �  �La8i�[�٬zF+�  �g�h�k<��@8K�  H���g�}7�ڒ�%�  ��g�mg�1&�3�   {4Wf����I�8�  �e�}�O���A�  8ӌ�d��_\���M�  P�4.d�ó�6D�  @��uc����2�I�  ��{�b��T�W�B�  `b��.�r�}�  X]�La��6MŞr<�  ��P�`���;ƥI�  p�η_��v�<�-�  �U�F^������9M�  ��\����̢N�  ��3e[��ݻ�k>?�   #J�Y�&�-D�  P�Z�X�m��4�I@�  @7eW��O���/�  �j�U���I�l�N�  �Ai0T��Wq�uI�  ��b�R��|m�:K�  �@VNQ�?|G¾d0�  `7��O�8��4�� �  �fX�L��z��B7C�  ��I�p4"%��H�  `/�G��:�
�WI�  `ȃ1D�/��!H�  @�%OA���A�9"I�  ��x�<�u*�6"dм  �7�xG��@�  @��O1���O(�;>�  ��'��8R�ؔN�   ;��*�2]��                   @G�?   �E�?   @D�?    C�?   �A�?    @�?   �>�?   @=�?   �;�?   @:�?   �8�?   �7�?    6�?   �4�?    3�?   �1�?   @0�?   �.�?   @-�?   �+�?   �*�?    )�?   �'�?    &�?   �$�?   @#�?   �!�?   @ �?   ��?   ��?    �?   ��?    �?   ��?   @�?   ��?   @�?   ��?   ��?    �?   ��?    �?   �
�?   @	�?   ��?   @�?    �?   ��?    �?   � �?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?    ��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   @��?    ��?   ���?    ��?   ���?   @��?   ���?   @��?   ���?   ���?    ��?   ���?    ��?   ���?   ���?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?    ��?   @��?   ���?   ���?    ��?   @��?   ���?   ���?    ��?   ���?   ���?    ��?   @��?   ��?   �~�?    ~�?   @}�?   �|�?    |�?   @{�?   �z�?   �y�?    y�?   @x�?   �w�?   �v�?   @v�?   �u�?   �t�?    t�?   @s�?   �r�?   �q�?    q�?   @p�?   �o�?    o�?   @n�?   �m�?   �l�?    l�?   @k�?   �j�?    j�?   @i�?   �h�?   �g�?    g�?   @f�?   �e�?   �d�?    d�?   �c�?   �b�?    b�?   @a�?   �`�?   �_�?    _�?   @^�?   �]�?    ]�?   @\�?   �[�?   �Z�?    Z�?   @Y�?   �X�?   �W�?    W�?   �V�?   �U�?    U�?   @T�?   �S�?   �R�?    R�?   @Q�?   �P�?    P�?   @O�?   �N�?   �M�?    M�?   @L�?   �K�?   �J�?   @J�?   �I�?   �H�?    H�?   @G�?                           �  �>Y� �"G=   � �>.ܶlW�E=   � �>jۋ�bH=     �>��^IL#=   � �>��(i�&I=   h��>g�ݟP'E=   p �>��*)��D=   � �>�&��N=   x �>.;ĝ��@=   H	 �>Qy�u�3=   �
��>�c���-=   �@�>R�ݡ�:==   ���>	��{M=    	@�>�����C=   `
��>b��ߔB=   � �>�td�C=   $��>���9��O=   � �>B� N��C=   ���>�j�&��==   ��>���.�<=    @�>`l�r�G=   ��>!���ls1=   � ?��8��=   �@?� �mN=   & ?��Ut�Q$=   X�?PiB�{^C=   ��?Gv�7��2=   �@?q�l��m+=   �?!�.j7�/=   d�?�L ��C=   �`?�m���	+=   P ?5Od%�	=   ��?�r����<   (�?*�Hga�2=   �@	?�C���I=   r 
?��s���A=   *�
?�GTi�A=   � `?�K�Ջ�D=   r" ?�Dp�`q=   L$�?��~���G=   4&�?����D=   �'@?�����E=   �) ?'P���<   �+�?f�4±cC=   �@?qW�n{;=   ��?�gC �i8=   ��?X�K�D=   P?G;��R"=   7�?�8΁3<L=   a?�rF҈K=   ^`?�_U�N=   ��?�;T��6=   � ?Ԛ����<   !�?q�W*#M=   ""�?�j�
�\M=   p#0?|I7Z#�/=   �$�?^��aDJ=   &�?��>,'1D=   B'@?�:�+NB=   �(�?�1z��@J=   * ?������3=   �+`?w�U4?�=   �,�?D��O=   ;.?$�b�� =   �/p?g)([|X>=   H1�?�>gV��=   �20?O�B��O=   *4�?bP�A��<   �5�?��e��4=   f7@?|[{�~*L=   9�?���ٹE=   t:�?G]����C=   '<P?�{m�u!K=   �=�?�
v\��4=   �??�����n=   fAp?�{7�!�O=   �B�?����=   �D ?�=u� �<=   �F�?�i&��-=   lH�?��o���N=   �I0?IT$7�QN=   �K�?Н��\�0=   �M�?0tЗ�I=   �OP?
�'��C=   uQ�?��4%@�@=   vS ?*�
qw�G=   ~U`?K ᴽ+=   �W�?F�Pn;�M=  ��, ?�]���K=  ��-8 ?�ƎI��M=  ��.h ?�5�m�3=   �/� ?�� ��M=   �0� ?�����I=   �1� ?�"���I=   �2 !?��y�$=  �4P!?�_	�D=  �.5�!?]��u�E:=  �"6�!?l�#�5=   J7�!?,����A=   u8"?��!y##�<  ��98"?�x�y�F=  ��:h"?bCڝ�D=   �;�"?u��RF=   =�"?2���w}=  �D>�"?�@(�6F=  ��? #?�'���A=   �@H#?43��A=  ��Ax#?uN}*�J=  �C�#?)�r7Yr7=  �]D�#?�.K="=   rE $?���r�=  ��F0$?3=1�Z1=   H`$?h|��=G=   gI�$?��ܩN�:=   �J�$?�4e��6=   �K�$?��{�<�9=  �=M%?uY�Pw�H=  ��NH%?��-*�8=  �Px%?�y�F�.=  �-Q�%?\9�;,=   �R�%?2�9Z�d@=   T &?~YK|=  �sU0&?WĻ��(J=  ��VX&?�R��IG=   X�&?W�	N=   �Y�&?�g�'9=   [�&?D�"^=   ���2)��$�   ����7�b�m�L�   Mӿ������(�   	ԏ��S��4�   ��_��	>��L�   |�/�����dM�   4���g±�8�   ����2�qڜ1�   �ן�qa�P�C�   Q�o�� ��%;9�   �?��_�0�C�   w��4g%6�L�   &���M��;k�@�   �ڿ�8�1�A�B�   ۏ�1�uB��   )�_����Y���   ��/�󓎣,:�   x����.Ճ^�-�   ������?�   �ޯ���ԝ�I�   -���:]=O>�   ��O�#w_jُB�   n�����(+E �   ���-�V~|_�   ����B}�_A�   C��K!ܨ�Y:�   ��_�5��G�   t�/��C���$>�   �����#���H�   m����-�
��M�   ���V���n@�   ���QU^�tA�   $�O��Ä�   ���þ��i�M�   @���K�8�|;2�   ���@�(�A�   V�����64�   ��o��ꬠTC�   9�?�&u����.�   ���~F�s:4�   �Կ��	��J�   ��_���L�II�   ����=�@�0(�   �ן��$�.�G��   ��?�}�3Rʏ3�   ����!|.4���   *ڟ�඄}��3�   �?�G"jm
>;�   ����*����O�   ���0 �:�O�   ������2K�;�   �޿�Q`���4�   ��_�� �ZD�   ���
���6�9�   *�
�����F�   �_
�T3ʢ�K�   ���	��M.�֢>�   ��	�@��_��@�   ��?	�1�\hU�   X������p�M�   &����J��x3�   ����Ҭ���   ���x�/h7�   8��L��v]E�   ����V���3�   ����B�v9�   r�_��c���M�   *����5&�L�   ���q����3�   ��?�:�R��$�   @���܎�$=�   ���K���'�   \�?��Ъ{�b>�   �����$E�vC�   ���I�w8�R'�   F��G�_j�,)�   ����+j�B�D�   |�_�`k�A�   ���%'r�BL�   ���	�T��E�   �_���GO�   ��� ��#i��#�    �� �;��^طH�   ��? �6(`J��J�   \����HB�5�   `����`��.11�   \�?��Q���D�   T����<VD��=�   D���Mϲk:UG�   ��?���,'��   �����h���UF�   ����U���ȘI�   �����t��@�5�   X�?��󕕠�4�   $������c��G�   ����y��/�C�   ������t�TM�   h�?���A�)E�   �����z�cϨN�   �����{���-��   <�?��G�#�?F�   ���}-w��F�   ����w���j'�   ���Q�x��   ��?����*
<�   4����	�,�   p��~ܾUY =�   �����˚�G�   ��쾂���p�7�   ���m�8�1<�   ����'����mN�   ��辙����L�   h���K��Y0�2�    ��̟q����   ���㾭v�Bfe9�   0���%��2�F�   ���ΥE��8�   ���߾�`�=�?�   ���ܾ��E=|
�   ���پu�M���   @��־��9��>�   ���Ӿ���9�6�   ���оk<
�xE�    ��˾�CqTR;�   ���Ǿ����dG�    �����G��gL�   @����_h�%?�   ������SS�@�                ��b��?�Wd���y>c��*GP��AiFC.ֿ      �?        53��=�?�͸�)a�<a�w>�,�?][S��q��n�C�?n�w���t�ӰY�?e�u��s�<���)kp�?&<��ߑ��țuE��?���K��a<����>��?5a1xH�<��lX��?
a�J.��<�Gr+���?qO���<���2���?R{�':@<���f��?{�N��k�Q[��?9�D9Ŗ��1l��*�?ǥl��Q��-���B�?�6�/��Q��ȘZ�?	��j@�<{Q}<�r�?u�׹A���ꍌ8���?k��#��u�o�[��?�hI{L[�<�\���?�.5�S����h1���?<d� n�<��"P��?��{�ߑ�֌b�;�?��J�uǍ<��}�I�?��~��<8bunz8�?rǶ~��<?��O�Q�?����U��<�|�eEk�?��@�3��<�c��߄�?}?�:L��������?U����<������?�8��
A�䦅��?�A�TG�<V/>����?�#�E�q<�1
��?�1�j�<1�L�p!�?|�眊<�d�<�?�Y6�!'�<�_�V�?(FN\�\��˩:7�q�?��B��:��f�m���?��<�������4ۧ�?��a�6�u���-��?�)]7����"4L���?���	ڊ<��E��?��V�#З�*.�!
�?x�0i�^���P��1�?�y_��ǁ�-�a`N�?π�z�H<W �Aj�?v�d�K��<�<�����?�b����s<����*��?V���b˙<'*6�ڿ�?�B쯗C}<������?3xj���<�,�v���?�WY�	���BfϢ��?i�v���O�V+4�?�<��z���]ʤQ�?����h���'�6Go�?��,��<�Ǘ���?��[ᕂ<)TH���?�GFL2�<�FY�&��?��i�K<<H!�o��?]�0���<	�v���?G�V�B⓼�U:�~$�?��@~���� ��4FC�?2��u<H��%"U�8b�?3Y�	���s�L�U��?d>�D�8`<�;f���?Ud�4ݛ���u��?�gV�r�/e<���?��<h:�k���Q�}��?��%<��t_��u�?�z��Gn��t��H�?�?;�el٨���gBV�_�?�m1WY$��?]�Oi��?,
�f�<��s��?/��w��2�0���?�M�L�<bN�6���?~y�]p<>T'�?*�mb�|���L��%�?�2�L����#FG�?��A��ֈ��D��h�?��ԛ�Ɵ��f��Ǌ�?:�|��<۠*B��?&K�V��<�D�2��?���2^�p�6w����?l��̅<���[�?#%X.y֝���Ͱ77�?�~���_g�R��DZ�?9�|Kv�PNޟ�}�?Ѕ|[����p��?2�Α�s���𣂑��?��q�F||<##�c��?nL�x�$x<e�]{f�?2�]IY��3-J�0�?�6�}\0�<]%>�U�?�A��n/��X�0�y�?�c��~˛<��yUk��?1�����<z�ӿk��?�l��4�����Z����?��]4͡�<f��)�?$�L�ޛ��O��3�?ׄ0^�b�:Y�rY�?�m���q��G^��v�?:�T~OXu�J�0���?.)T������K���?��-z�=�<	�[���?r�k?�����R�ݛ�?�HP�e�<z��_�@�?
ƃ�7E�<K�W.�g�?�<H�M��<���m��?D\�H��q<i��� ��?�I���u<��]U��?r��S;؍�|�J-�?�zyC7�����/�?w��q{H������X�?7[��<�����?�������2���?2�mi #�<`��!��?��xWڒ<_�{3���?[KOͥ��)��F&�?�z�'����?��.P�?�̩����<�L��Qz�?��"Ւ<ڐ�����?�(�#����g�-H��?���󓜼'Za���?�����ǝ<��k7+%�?C�����<@En[vP�?���-�ә<����{�?	5����ؐ�����?���SH�<�q�+���?�ye�t�b<      8C      8C������ ������       �?      �?��������������1g���U?���k�?wN�o���?�ł����?�9��B.�?   �����   @G��     �      �      ��       �      ��      �             ��        ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx                            8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?       �           �����   �����    ���UUUUUU�?333333�?�m۶mۦ?颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?       �9��B.�@  ׽2b      �              8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?\3&���-DT�!	�\3&��<-DT�!	@       �           �����   �����    ���                UUUUUUſ333333���m۶mۦ�颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?      �?       �9��B.�@  ׽2b      �              �7                              �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������                                      �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      �      �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow       �      ���������������-DT�!�?-DT�!��RUUUUU�?        v�F�$I�?������ɿ��3Y�E�?#Y��q���n����?��;
9��� ��/I�?hK����d��?81�U����H!G�?��#�$�����0|f?�K�RVn���TUUUU�?        ~I�$I�?g����ɿHB�;E�?����q���{雮?�x��֚��                   �      �?       @       @      �?      �?      @>��1|�MC              ������ ������ ������B������B  �����  ����� 8��B.�?0gǓW�.=        ����������������              �?      �?                      0C      0C      ��      �     �     �U�	�I�? ���Ͽu}�M�Uſ�UUUUU�?Sz�����?     �      �?      �?     ��?     ��?     �?     �?     ��?     ��?     �?     �?     ��?     ��?     B�?     B�?     ��?     ��?     r�?     r�?     �?     �?     ��?     ��?     N�?     N�?     ��?     ��?     ��?     ��?     B�?     B�?     ��?     ��?     ��?     ��?     H�?     H�?     ��?     ��?     ��?     ��?     b�?     b�?     �?     �?     ��?     ��?     ��?     ��?     F�?     F�?     �?     �?     ��?     ��?     ��?     ��?     B�?     B�?     �?     �?     ��?     ��?     ��?     ��?     V�?     V�?     �?     �?     ��?     ��?     ��?     ��?     z�?     z�?     F�?     F�?     �?     �?     ��?     ��?     ��?     ��?     ��?     ��?     R�?     R�?     $�?     $�?     ��?     ��?     ��?     ��?     ��?     ��?     t�?     t�?     J�?     J�?      �?      �?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     \�?     \�?     6�?     6�?     �?     �?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     ��?     b�?     b�?     B�?     B�?      �?      �?      �?      �?                  <����?N~�'��<  x�z�?��'�*$=  �#�f�?�$/��= @�0�?@A�S��1= �c�E�?�Pa�B== `�R�?Dj0Q:W$= ��>m��?��Lyc>= �*p%�?���?C;0= ��|���?�Ix�"�<= ``ә�?��y M== �or�O�?��+C��== ��v��?�����R1= PQ	��?��Ӏb= @��P�?�5M[g?= �V���?d+��[7= ������?n��B�>=  kz�*�?�w�#8= 0�nط�?C�#�7= �{���?Di�00= �ˮf�?�j -= x���)�?���}z�=  ����?��0$= H�V��?����o�= X��a�?��;�M_8= @��?�����5= ����?�^���@'= �L$��?��/r(= � <�?�vT�� 3= ��?���?��Cg��?= 0��Ә�?W/f�1= `(J�?Dk����0= h��#��?@� �6= �۫���?��_��= �|�D�?�&�?4j<= '����?Q���n�&= �ַ��?�l����= �Ð6�?�DX�,4= �����?��-Q�2= �xb�t�?�W��E��< �.l�?��7�w�,= ���Ȭ�?l�>= �ɥ�%�?��Nl,"= �@\r�?�?� t�8= 85�R��?ӇӜ��= L.��	�?�>)g�= Ը�3U�?�Ӱ��== �����?h���Xg+= �og���?�����X= ��ذ0�?{fHn�= <��w�?y�5s3R6= ��)��?��a8��< O4W�?4�bV�0= ����L�?�4���@= ���@��?�X��ۓ4= Tk���?>�_��(=  ����?�*��o= �@�[c�?�����,= $4b��?d����O"= lx���?#60���8= ě&m*�?ɉ�h"0= �בl�?�n6ѯ{�< 9[P��?�ce�zb�< $����?�F�8"= 8��B.�?0gǓW�.=�������             ��      �@      �        	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ =                      �       �      ��      ������    ����    ��      ��            8C      8C      0<      0<��+eGW@��+eGW@  ��B.�?  ��B.�?:;����=:;����=�ѱt�?Z�fUUU�?���&WU�?{������?                Mu�{�<`�w>�,  �g5RҌ<t�ӰY  a��aN�`<țuE�  l{�]���<��lX�  ќ/p=�><���2��  ؼcnQ�<P[� {8�&TŤ<�-���B �?RbSQ�<zQ}<�r �S?���<u�o�[� _/:>��<��h1�� �æDAo�<֌b�; �������<8bunz8 ���+G�<�|�eEk 1�	m���<����� �
r�7�<䦅� ���MuM�<�1
� J��]9ݏ<�d�< )}̌/�<ʩ:7�q �^�s)ҧ<���4ۧ mL*�H��<"4L�� ��%F��<).�!
 ��`�cC<-�a`N y����n<�<���� ��z�ΐv<'*6�ڿ 	*(�̃�<�,�v�� ���	�<�O�V+4 ���5�<�'�6Go 	T��c�<)TH�� 5�d+�2�<H!�o� 
���<�U:�~$ �s ��<$"U�8b qU�M��<�;f�� �GΆ�+�<.e<�� �o � �<s_��u ���"a�<�gBV�_ ��F�D�<��s� Ul֫��e<bN�6�� �g�����<�L��% ���<�D��h ����/��<۠*B� D_�Y��{<6w��� <(��`�<��Ͱ77	 �b� ��<ONޟ�}	 'Α+��q<�𣂑�	 �.�X4m�<d�]{f
 ����|'�<\%>�U
 �Zsn�i�<��yUk�
 �3˒w�<��Z���
 �-�f$�<�O��3 ���.�<F^��v ��_
��t<��K�� ��0�ns<�R�ݛ �Y	я��<K�W.�g h�l,kg<i��� � ���6	p�<{�J- �=���t<����X ����PZ�<�2�� ��Js��<^�{3�� ӈ:`�t<�?��.P &I	�'o�<ِ����  �A�Î<'Za�� ��1�d�<@En[vP �͑M;�w<ؐ����       �?       �9��B.�@  ׽2b      �        �������         0<  0<�dW�dW                �,��d�?                        =��U�&�?UUUUUU�?                �}=mm?�?                �u+E6�W?�����?                      �?                        �_CN�?�?        F�n<�t�?        u[�c��?�#�Xu�?�7�&�?�I�v�*�?��w�|u?!u$�8�?"Y�Nu?-HF���?0[��d? cf>	�?����c?����?�-[��6�?���N}X<      �?�]���݃?                ��'Z4�?        �e-CS�?        F���?��,��w�?(F_�e��?�X2CQ��?	ُ�㈏?�wT��?�/V�W��?#�(�7�?��� L�?�hC!�߶?c�(��y?�-�˶?X1U��u�?�?Y��.<      �?P��B�?                >S�Ŏ�?        �6�	�Ӷ?        �'��P9�?��z�^3�?��
΂��?&1yA��?�(+_�R�?m�Y��?�}�"��?�Ɵ�lW�?P),��H�?,��b��?�����?@��?��?�c\5j�?=��Mpm�      �?c��+���?                Bp�VV��?        Q9V�%�?        ]|=3�?.����?|��_P��?�%�����?ػZq\�? ,6���?�5DKBӹ?�@IK��?�Xf���?v������?�'���?+�3���?2���y��?g��/�p<      �?7C���?                ����?        E�D;��?        ��h7�r�?��=���?(��r�?�EV�w�?��У��?�����?0�SM`��? ��?3��?/��*2�?5�6Y�z�?�Ʊ���?�G�e�?�4��?�%��KV��      �?�r��H�?                �I,+���?        ��U&X>�?        �i�.��?�c4���?����?�����?��N�T�?��j8�6�?�f*"!��?~w�"�?nJ�R��?1 ��7!�?|�GD|�?���?���*�a�?�}� Ũ�<      �?ƼpAؒ�?                ZM��$^@        ]�>�=�@        Z��7@�abK���?؝Z��@ �t���?��,��@�T��4s�?�ag�@Xp�M� @�D�$_�@�n}in @��)�M�@֐��@P(�* C�?� ��mz�       @�E3�&�Կ                fY�eY�!@        �,��d&@        #7̓B�,@       @=��U�&2@UUUUUU@9E4�7@������
@�}=m=@@ 8�λB@[�[�@�u+E6�G@����@      �?               @                        ӸHO��3�        oX�� ?        �%��
���#�Z��."S-�>Q�!�r�?�M%���ᾎ;���Ǆ�c�d3�>����$9t?��Jy��������A]�VJ��]�>Q��䫢I? ��Z�Iο7t�`�=        �cH���?      �?    ������ZS �+�        ߏ�?        ��Y�9�m|1�~��-g���>b/[E�?8��QSվ��7��K�����Ǔ��>���p?[j3�H��X�&
C�U��x����>Xzv�C?  �*�ɿa�#wi#:�        ��w�B��?      �?    �������x#�        �qQ���?        �Ly�a���F������5d����>2�*�q�?����ɾ���?c3y��Ɵ0��>q澺�k?��������g\>{�O�>>��u��>�����=? ��)�IſX��3{9�        l���f�?      �?    ����V��}X9�        ܈��?        +*tsJ�E�X*��y�hU&��>��3��H�?��ܨ9�����ԪF�r�������>�)��(�g?����V����t��F�cf���y>?���p�6? �������K�=��3�        il���?      �?    �����Kk�        0vB-�G?        � 8��d��l������M���V�>|s`���?���P���t��"�!k���?J�I�>΃+�תd?�s{c|H��Y"��?���X��:n>�/��/�2? �6�G�������^�        #���f��?      �?    ����d�čD�        o=���z�>        -�B���վ��y%�#����(A�>ō�:��?S��/�|��o3fW�|a��D	`�N�>���F�b?���k��t�	L�R�3�e����c>D���f�/? @��b̰��k���        �ع��?      �?    �����"�]�)��        E��}��>        ��r>ľ>�n���z�ru���>�Cԑ��?lf6	n����oP�"Q�?�m˹A�>���fǰa?+�kW�Zb����I#�݄,[>�=�h��,? ��nĠ���}�P=        �Ȣ��_�?      �?    ����                ��+�j�>                        &D�(�>l�l��?                b��Ĳm�>g�jVa?                \�yN�W>�4�w�+?                        UUUUUU�?      �?    �����"�]�)�>        E��}��>        ��r>�>>�n���z?ru���>�Cԑ��?lf6	n�>��oP�"Q??�m˹A�>���fǰa?+�kW�Zb>���I#?݄,[>�=�h��,? ��nĠ?��}�P�        �Ȣ��_�?      �?    ����d�čD?        o=���z�>        -�B����>��y%�#�?��(A�>ō�:��?S��/�|�>o3fW�|a?�D	`�N�>���F�b?���k��t>	L�R�3?e����c>D���f�/? @��b̰?�k��=        �ع��?      �?    �����Kk?        0vB-�G?        � 8��d�>�l����?�M���V�>|s`���?���P��>t��"�!k?��?J�I�>΃+�תd?�s{c|H�>Y"��??��X��:n>�/��/�2? �6�G�?�����^=        #���f��?      �?    ����V��}X9?        ܈��?        +*tsJ�>�E�X*�?y�hU&��>��3��H�?��ܨ9��>��ԪF�r?������>�)��(�g?����V��>�t��F?cf���y>?���p�6? �����?�K�=��3=        il���?      �?    �������x#?        �qQ���?        �Ly�a�>�F����?�5d����>2�*�q�?�����>���?c3y?�Ɵ0��>q澺�k?������>�g\>{�O?>>��u��>�����=? ��)�I�?X��3{9=        l���f�?      �?    ������ZS �+?        ߏ�?        ��Y�9?m|1�~�?-g���>b/[E�?8��QS�>��7��K�?���Ǔ��>���p?[j3�H�>X�&
C�U?�x����>Xzv�C?  �*��?a�#wi#:=        ��w�B��?      �?    ����ӸHO��3?        oX�� ?        �%��
?��#�Z�?."S-�>Q�!�r�?�M%����>�;���Ǆ?c�d3�>����$9t?��Jy���>����A]?VJ��]�>Q��䫢I? ��Z�I�?7t�`��        �cH���?      �?    ����fY�eY�!�        �,��d&@        #7̓B�,�       �=��U�&2@UUUUUU@9E4�7�������
��}=m=@@ 8�λB�[�[���u+E6�G@����@      �               @                        ZM��$^�        ]�>�=�@        Z��7��abK����؝Z��@ �t���?��,����T��4s���ag�@Xp�M� @�D�$_���n}in ���)�M�@֐��@P(�* C�� ��mz<       @�E3�&�Կ                �I,+���        ��U&X>�?        �i�.��c4�����?�����?��N�T����j8�6��f*"!��?~w�"�?nJ�R���1 ��7!�|�GD|�?���?���*�a��}� Ũ��      �?ƼpAؒ�?                ���߿        E�D;��?        ��h7�rۿ��=���(��r�?�EV�w�?��У�׿�����0�SM`��? ��?3��?/��*2Կ5�6Y�z⿛Ʊ���?�G�e�?�4���%��KV�<      �?�r��H�?                Bp�VV�̿        Q9V�%�?        ]|=3ſ.���߿|��_P��?�%�����?ػZq\�� ,6��ڿ�5DKBӹ?�@IK��?�Xf��䵿v�����ӿ�'���?+�3���?2���y�ڿg��/�p�      �?7C���?                >S�Ŏ��        �6�	�Ӷ?        �'��P9����z�^3տ��
΂��?&1yA��?�(+_�R��m�Y�п�}�"��?�Ɵ�lW�?P),��H��,��b�ſ�����?@��?��?�c\5jӿ=��Mpm<      �?c��+���?                ��'Z4��        �e-CS�?        F������,��wʿ(F_�e��?�X2CQ��?	ُ�㈏��wT�¿�/V�W��?#�(�7�?��� L��hC!�߶�c�(��y?�-�˶?X1U��uɿ�?Y��.�      �?P��B�?                �_CN�?��        F�n<�t�?        u[�c����#�Xu���7�&�?�I�v�*�?��w�|u�!u$�8��"Y�Nu?-HF���?0[��d� cf>	棿����c?����?�-[��6�����N}X�      �?�]���݃?                ���m0_$@���m0_$@      xC      8C @DT�!�?  DT�!�? @gg��2�  LL#�F=J47ࢨ:Esp.��:�3gg��2=      �?  ������               �      `C      �<      �<      �        c c s =     U T F - 8   U T F - 1 6 L E     U N I C O D E   ccs=    UTF-8   UTF-16LE    UNICODE _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh            ������ ������      ��?     ��?������B������B   ����   ���� x�PD�?X�1�=        ����������������              �?      �?                      0C      0C      ��      �     �     ��Η��5@=�)d	��U�5j��%��5��j�?��~��@5�w��z�A.�lzZ?                          �
�|?�Q-8>=  ޶�W�?0��	k8= ��ޮp�?�x�9=  >�.ښ?pn��5= �Y�ح�?�  	Q*=  c����??���b6= ��Y�?�T�?�=  ��>�?����W�!= @�-32�?D���z= ��p(�?vP�(��= `����?�US?�>= �e��?�g���7= `ŀ'��?�bͬ�/= ��^s�?�}�#��= �J�wk�?zn��= ��Nָ?�LN�� 9= @$"�3�?5Wg4p�6= ��T���?�Nv$^)= ��&�?��.�)��< �l��B�?�M���%= `j���?�w����*=  <śm�?E��2=  ެ>�?����E�= �t?��?����= �O�Q�?�w(@	��< ��0��?Ac��0= Pyp��?dry?�= ��St)�?4K��	�>= ���$��?Qh�BC .= 0	ub�?-����0=  ���?a>-�?=  ����?Й��,��<  (lX �?�T@b� == P����?�3�h,%= ��f�?�?�#���� = �V��?ߠϡ��6= ����Y�?���z $= ��G��? $�l35= @��n�?[+���3= �Rŷ �?s�dLi�== p�|��?r�x"#�2= @.���?|�U��2=  lԝ��?r��F�= �a��?����4= ��Y��?sl׼#{ = `~R=�?�.�i�1= ��,��?���� = ��vX�? ���= p����?h���}s"= �	E[
�?%S#[k= ��7�H�?����j= �!V1��?��}�a2= �jq��?2�0�J�5= ������?����5= x¾/@�?��"B <1= �i�z�?�\-!y�!= X�0z��?~��b>�== �:���?�#.X'= HBO&�?��(~= x�bb�?.�= �C�q��?y7��i9+= �v���?����:= 0����?2ض��8= x�PD�?X�1�=     ��?     ��?     Q�?     Q�?    ���?    ���?    ���?    ���?    ��?    ��?    ���?    ���?    �]�?    �]�?    P�?    P�?     ��?     ��?    �U�?    �U�?    (��?    (��?    `��?    `��?    �_�?    �_�?    ��?    ��?    ���?    ���?    �z�?    �z�?    �1�?    �1�?    p��?    p��?    ��?    ��?    (e�?    (e�?    @#�?    @#�?    ���?    ���?    `��?    `��?    hk�?    hk�?    �,�?    �,�?    x��?    x��?    ���?    ���?     ��?     ��?    �N�?    �N�?    x�?    x�?    p��?    p��?    ��?    ��?    �~�?    �~�?    HN�?    HN�?    ��?    ��?    ���?    ���?    ���?    ���?    p��?    p��?    Xi�?    Xi�?    �?�?    �?�?    ��?    ��?     ��?     ��?    ���?    ���?    8��?    8��?    s�?    s�?    pI�?    pI�?    �&�?    �&�?    � �?    � �?    ��?    ��?    �o�?    �o�?     *�?     *�?    ���?    ���?    `��?    `��?     Z�?     Z�?    ��?    ��?    0��?    0��?    ���?    ���?    PY�?    PY�?    ��?    ��?    `��?    `��?    ��?    ��?    pm�?    pm�?     /�?     /�?    ���?    ���?     ��?     ��?InitializeCriticalSectionAndSpinCount   kernel32.dll     Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ()  >=  <=  /   ->* &   --  ++  *   ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        x�p�d�X�L�@�4�,� ��k4t�X�D�$���� h �����������ܒؒԒВ���#̒ȒĒ�#�'���'��K���-����������������������������t�h�`�T�<�0����ܑ����|�X�<����А����������d�\�P�@�$��܏����`�D� ���Ў����k4GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL  ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp              �U��?�wB%�K�=      �?   �[��?(�6N�g�=      �?   $�?V�`t� >      �?   ��տ?��2n{a>      �?   ����?��M��=      �?   H{��?{4�r>      �?   Pא�?"�"�>      �?   �u[�?��*��>      �?   ����?G�0��_(>      �?   4wb�?��i^^?(>      �?   ��0�?p3���>      �?   @��?F��M>      �?   8M��?�B�V��>      �?   ��d�?}B��a.>      �?   ȴ�?d�����>      �?   g��?�ߊ��>      �?   �@�?�f\���*>      �?   �~e�?�-��f>      �?   �]%�?D	�G��?>      �?   ���?�\����>>      �?   X���?�1��#>      �?   �E�?��h��>      �?   �?��?�ⳇ��>      �?   ����?�$	�49>      �?   x�8�?k���0H<>      �?   ����?r��ش8>      �?   8fm�?�"m>">      �?   ħ �?[��<c�'>      �?   �k��?"���%>      �?   ���?݉@fR�8>      �?   ����?��T���:>      �?   T�!�?3&�F>      �?   � ��?<����[#>     ��?   �%�?�Y:/(A6>      �?   ����?��N��2>     ��?   8O�?�r�!'	>      �?   ��r�?���8{K>     ��?   �p��?9��l�9$>      �?   �
G�?�aj	�i9>     ��?   T|��?'\�|#<>      �?   $��?�}�dj�#>     ��?   �Wn�?׈MVx:>      �?   ,���?1�8o,>     ��?   D�$�?	c�/�
>      �?   @ |�?��x7|�1>     ��?   |���?��9>      �?   p #�?�IA��u=>     ��?   �s�?�x ٴ4>      �?   p���?edf�&�.>     ��?   ,�?��f���A>      �?   h�*�?v����2>     ��?   $gN�?RE\��K>      �?   �q�?'^��IE>     ��?   DΒ�?��&a��H>      �?   L���?�&KrQF>     ��?   ,���?�#/�'�>      �?   إ��?]X�c�?>     ��?    ��?�Ԯ}�>      �?   �e.�?�IdW�A>     ��?   �K�?���ΐ?>      �?   Xg�?��4*�A>     ��?   _��?�[�ǆJ>      �?   ���?1���0H>     ��?   ���?�hc#�]G>       @   ,*��?�Q�x
�F>     @ @   p���?ek�R�.N>     � @   �� �?�Ӿ�n@>     � @   �b�?�����O>      @   $Q/�?CJ���O>     @@   ��E�?������G>     �@   �[�?�3E�{A>     �@   T�p�?�SfI�S:>      @   X΅�?B6)�1�<>     @@   �3��?>ځ���7>     �@   $��?s(��N>     �@   @���?V�
6�f=>      @   (���?��{��>     @@   (W��?��-�Jg >     �@   ����?��"a�PK>     �@   xm�?,S��ڤ6>      @   ���?�6��hb">     @@    �-�?�k,�<>     �@   X�>�?�0����=>     �@   �O�?�׀IX�H>      @   �-_�?���
@>     @@   ��n�?���2E>     �@   �P~�?�=�ő�8>     �@   lj��?�[j&,>      @   L7��?��x��82>     @@   ����?c�#V�B>     �@   0��?7ڨ.�Y>     �@   P���?�[�p&>      @   ؔ��?h4�M��A>     @@   � ��?E�p�l E>     �@   �+��?�o�$�E>     �@   h��?\���*�K>      @   ���?-�?��B>     @@   P8�?�(l�|�@>     �@   �p!�?u���@�J>     �@   @p-�?�V��1>      	@   �89�?����5>     @	@   <�D�?��ƀ�7>     �	@   h)P�?R`D�OG>     �	@   �T[�?9%� ��K>      
@   �Mf�?��/�<>     @
@   �q�?�Ò��?>     �
@   �{�?4��2G<>     �
@   L��?Â���|/>      @   �Y��?���s�
@>     @@   �k��?��Ò�a@>     �@   XS��?x(3��u8>     �@   ���?v�O,ib>      @   ȥ��?�&L͒C>     @@   ���?��}��L>     �@   �X��?Lo����>     �@   �x��?-�Ϡ�9>      @   �s��?6FID?9>     @@   8J��?����gsL>     �@   d���?��y>     �@   ���?>�&�09C>      @   ����?
��<�A>     @@   (J�?I�V	C>     �@   `w�?��^@�N>     �@   ���?�#��%�@>      @   �s�? �M�K>     @@    D'�?ή�Q��->     �@   ��.�?9!���G>     �@   ��6�?.����1>      @   >�?.1�NcB>      @   �cE�?�sǔ�1>     @@   L�L�?�n�HN>     `@   H�S�?�W��$>     �@   8�Z�?
Ȃ�q�;>     �@   ��a�?N�/�[7>     �@   (�h�?�=�mC>     �@   0oo�?�H75M>      @   Hv�?P��.�#>      @   �|�?�G���7>     @@   �*��?�#4��2I>     `@   ����?o���oJ>     �@   ����?���-��#>     �@   ���?�h��%F>     �@   @��?R�x^D>     �@   PP��?�� s�@>      @   4L��?P�_!
�#>      @   4��?��:#�G>     @@   L��?qg�:&J>     `@   Hɹ�?5L$.��4>     �@   \w��?!�1�C>     �@   ���?���[<>     �@   D���?��<���=     �@   ���?��
~���=      @   �y��?������B>      @   ����?�~.���4>     @@   h��?��u�|�8>     `@   �E��?A8yL;>     �@   �h��?��41��C>     �@   �{��?-���+oF>     �@   $��?x���O>     �@   s��?�՝m�T2>      @   �W��?����=>      @   �-�?î�\�=>     @@   ��?���\=�=     `@   ��?j\&">     �@   �X�?��1�D>>     �@   ���?�#O#`�I>     �@   ��?�}���0>     �@   ��?���F\IE>      @   t{#�?��ׯ,B>      @   0�'�?�E� ]�$>     @@   ,>,�?��ކ?5>     `@   ��0�?��iIqE>     �@   ��4�?�ha�;>     �@   �9�?��A���D>     �@   �.=�?̤KF�w�=     �@   DMA�?�����=      @   `E�?ap�I0�H>      @   �gI�?��:���->     @@   �cM�?��%Q>     `@   @UQ�?Ly5ښoE>     �@   �;U�?v�g�0�/>     �@   �Y�?jv�U�G>     �@   �\�?�����yK>     �@   ,�`�?A%My��>      @   md�?���H>      @    h�?�p���M>     @@   0�k�?k��}<>     `@   �ho�?����f7O>     �@   ��r�?���}�O>     �@    �v�?+��i�I>     �@   @z�?�b�B'=>>     �@   `�}�?Z����M>      @   ����?1�����M>      @   �a��?R�~���=     @@   t���?QNT	��B>     `@   x��?�W3c�L>     �@   g��?�+(����=     �@   D���?q���J�K>     �@   L��?� ;,*>     �@   8!��?������D>      @   ,O��?� ����E>      @   Du��?��in]D>     @@   ����?%����3F>     `@   P���?^��F"VM>     �@   ����?�}�30}->     �@   @���?�~F	y�;>     �@   ����?l	R(>     �@   躰�?��\�7`>      @    ���?�dg���;>      @   ���?�;Sv�@E>     @@   <|��?�����M>     `@   �Y��?|}�;�2>     �@   ,0��?�<v��G>     �@   $ ��?̯�/p�">     �@   ����?���\(0>     �@   |���?[s$���F>      @   I��?�d�ӔV>      @   T���?���0)LK>     @@   h���?�)�5G�5>     `@   XY��?�|��zJ>     �@   @���?W�޾�L?>     �@   0���?����6:>     �@   <3��?��Q���B>     �@   x���?7o��/�M>      @   �Q��?�Kc�Z�0>      @   ����?�z-�A5>     @@   Z��?"B�DcI>     `@   ����?��`I�.>     �@    L��?L�d�%>     �@   ���?"�l"w �=     �@   �(��?�?��!>     �@   ���?��j^�J>      @   8���? ϞH��0>      @   LL��?���%�C>     @@   T���?��J�+N>     `@   d���?;l�>�0>     �@   �B��?�^{v�@>     �@   Ȋ��?�@Y˕B>     �@   @� �?T�l���0>     �@   ��?w4n4>      @    G�?�oN�=�;>      @   h|�?�L�{�/>     @@   <�	�?B�nu5>     `@   ���?���`�,+>     �@   d�?����5>     �@   �$�?l��  >     �@   �C�?~+^��M>     �@   �^�?�PK�QD >      @   ,u�?^{�#tF>      @   |��?�^4K�� >     @@   ���?��4�O
>>     `@   ���?XEړ� J>     �@   ���?(�gԹ�,>     �@   �� �?43-spF>     �@   ��"�?P`E5�+*>     �@   ��$�?=�QQ�D>       @-DT�!�?\3&��<                                                                                                                                                                                                                                                                                  ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  Dec Nov Oct Sep Aug Jul Jun Apr Mar Feb Jan Sat Fri Thu Wed Tue Mon Sun SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    1#QNAN  1#INF   1#IND   1#SNAN  CONOUT$     H                                                             `�  RSDS~�����M�?�|�<Y\   C:\Program Files\MAXON\CINEMA 4D R12\plugins\rhinoio\obj\rhinoio_Win32_Release.pdb             ����ķ    �       ����    @   ��$�        ����    @   �           �ķ                <��           �,���ķ    <�       ����    @   �            h�\�           l�x���    h�       ����    @   \���        ����    @   ��           ����               ظ�ķ    ��       ����    @   ȸ            ���           $�,�    ��        ����    @   �            ��\�           l�t�    ��        ����    @   \�            ���           ����    �        ����    @   ��            0��           ���    0�        ����    @   �            \�4�           D�L�    \�        ����    @   4�           x����ķ    ��       ����    @   h�            ����           Ⱥܺ���ķ    ��       ����    @   ��            ���           �(���    ��       ����    @   �            ��X�           h�x�(���    ��       ����    @   X�           �����ķ    �       ����    @   ��            0��           ������ķ    0�       ����    @   �            P�8�           H�X�(���    P�       ����    @   8�            t���           ������    t�       ����    @   ����        ����    @   ܼ           ���                ���           � �    ��        ����    @   �            $��           `�h�    ��        ����    @   P�            ���           ����    �        ����    @   ��            4��           ���h�    4�       ����    @   �            d�,�           <�D�    d�        ����    @   ,�            |�t�           ����D�    |�       ����    @   t�            ����           оؾ    ��        ����    @   ��            ���           �$�D�    ��       ����    @   �            ��T�           d�t�$�D�    ��       ����    @   T�            ��ܼ            ���           ȿп    �        ����    @   ��            <� �           ��    <�        ����    @    �            X�H�           X�`�    X�        ����    @   H�            x���           ����h�    x�       ����    @   ��            ����           ����    ��        ����    @   ��            ��$�           4�<�    ��        ����    @   $�            ��l�           |���<�    ��       ����    @   l�            ���           ������<�    �       ����    @   ��@�       ����    @   �            ���<�                \�@�           P�X�    \�        ����    @   @�            ����           ������<�    ��       ����    @   ��            ����           ����    ��        ����    @   ��            �� �           0�<�<�    ��       ����    @    �            �l�           |���    �        ����    @   l�            <���           ����    <�        ����    @   ��            p���           ��    p�        ����    @   ��            ��D�           T�`�<�    ��       ����    @   D�            ����           �������<�    ��       ����    @   ����       ����    @   ��           �����<�    ��       ����    @   (�           8��<�                ����            ��l�           |���    ��        ����    @   l�            ���           ������    �       ����    @   ��            $� �           � ��<�    $�       ����    @    �            D�P�           `�p��<�    D�       ����    @   P�            d���           �����<�    d�       ����    @   ��            ����            ����<�    ��       ����    @   ��            ��@�           P�X�    ��        ����    @   @�            ����           ����    ��        ����    @   ��            ���           ����    �        ����    @   ��            0��           (�0�    0�        ����    @   �            h�`�           p�x�    h�        ����    @   `�            ����           ����    ��        ����    @   ��            ����            ��    ��        ����    @   ��            �8�           H�P�    �        ����    @   8�            8���           ����    8�        ����    @   ��            p���           ����    p�        ����    @   ��            ���            �(�    ��        ����    @   �            ��X�           h�p�    ��        ����    @   X�            ���           ����    �        ����    @   ��            8���           �����<�    8�       ����    @   ��            \�8�           H�X��<�    \�       ����    @   8�            t���           �����<�    t�       ����    @   ��            ����           ������<�    ��       ����    @   ��            ��(�           8�@�    ��        ����    @   (�            ��p�           ����    ��        ����    @   p�            ���           �����<�    �       ����    @   ��            @��           �(���<�    @�       ����    @   �            l�X�           h�|����<�    l�       ����    @   X���       ����    @   ��           �����<�                ����           �����<�    ��       ����    @   ��            ��8�           H�P�    ��        ����    @   8�            ���           ����    �        ����    @   ��            <���           ����    <�        ����    @   ��            l��            �(�    l�        ����    @   �            ��X�           h�p�    ��        ����    @   X�            ����           ����    ��        ����    @   ��            ����           �� �    ��        ����    @   ��            , 0�           @�H�    ,         ����    @   0�            \ x�           ����    \         ����    @   x�            � ��           ���� ��<�    �        ����    @   ���        ����    @   �           ,� ��<�                � P�           `�x������<�    �        ����    @   P��        ����    @   ��           �������<�                � ��           ��������<�    �        ����    @   ��            @�           P�`��<�           ����    @   @�            0��           ���������<�    0       ����    @   ��L       ����    @   ��            ������<�                l(�           8�D���    l       ����    @   (�            �t�           ����(�    �       ����    @   t�            ���           ������    �       ����    @   ��           ��p�    �       ����    @   ��           @�L� �    ,       ����    @   0�            \|�           ����D���    \       ����    @   |�            ���           ������(�    �       ����    @   ��            ��           ,�<��p�    �       ����    @   �            �l�           |�������    �       ����    @   l�            ���           ����L� �    �       ����    @   ��             �           �,��<�            ����    @   �            � �            p�           �����<�           ����    @   p�            0��           ����    0        ����    @   ��            `�           � �    `        ����    @   �            �P�           `�h�    �        ����    @   P�            ���           ����    �        ����    @   ��            ���           ����    �        ����    @   ��            4(�           8�@�    4        ����    @   (�            hp�           ����    h        ����    @   p�            ���           ����    �        ����    @   ��            � �           ��    �        ����    @    �             H�           X�`�             ����    @   H�            0��           ����    0        ����    @   ��            \��           ����    \        ����    @   ��            � �           0�8�    �        ����    @    �            �h�           x���    �        ����    @   h�            ���           ����    �        ����    @   ��            ��           ��            ����    @   ��            P@�           P�X�    P        ����    @   @�            ���           ����    �        ����    @   ��            ���           ����`�    �       ����    @   ��            ��           ,�8���    �       ����    @   �            h�           x�����           ����    @   h�            <��           ������    <       ����    @   ��            p �           ���    p       ����    @    �            �L�           \�h�8�    �       ����    @   L�            ���           ������    �       ����    @   ��            ���           �� ���    �       ����    @   ��            00�           @�L��    0       ����    @   0�            h|�           ����    h        ����    @   |�            ���           ����<�    �       ����    @   ��            ��            �,�<�    �       ����    @   �            �\�           l�t�    �        ����    @   \�            ���           ����t�    �       ����    @   ��             	��            ��<�     	       ����    @   ��            T	<�           L�\��<�    T	       ����    @   <�            p	��           ����    p	        ����    @   ��            �	��           ����    �	        ����    @   ��            �	�           ,�4�    �	        ����    @   �            
d�           t�|�    
        ����    @   d�            @
��           ����    @
        ����    @   ��            p
��           ��    p
        ����    @   ��            �
<�           L�X�(�    �
       ����    @   <�            �
��           ����,�    �
       ����    @   ��            �
��           ����p�    �
       ����    @   ��              �           0�<�X�            ����    @    �             l�           |�����            ����    @   l�            @��           ������    @       ����    @   ����        ����    M   (�            \ �           0�<�X�    \       ����    @    �P        ����    M   @�            |��           ������    |       ����    @   ��p
        ����    M   ��            ���            ����<�    �       ����    @   ��            �@�           P�X�    �        ����    @   @�             ��           ����             ����    @   ��             ��           ������            ����    @   ��            <�           ,�8���    <       ����    @   �            dh�           x���    d        ����    @   h�            ���           �������<�    �       ����    @   ��            ��           ��    �        ����    @   �            �L�           \�p����<�    �       ����    @   L�            ���           �������<�    �       ����    @   ��            ���           ���    �       ����    @   ��            @�           P�d����<�           ����    @   @�            4��           �����    4       ����    @   ��            X��           ������<�    X       ����    @   ��            @��            tH�           X�h���<�    t       ����    @   H�            ���           ������    �       ����    @   ��            ���           �� �<�    �       ����    @   ��            �0�           @�P���<�    �       ����    @   0�            ��           ������<�           ����    @   ��            $��           ������<�    $       ����    @   ��            L �           0�@���<�    L       ����    @    �            tp�           �����<�    t       ����    @   p�            ���           ������<�    �       ����    @   ��            ��            �0��<�    �       ����    @   �            �`�           p���0��<�    �       ����    @   `�            ���           ����0��<�    �       ����    @   ��             �           �,�0��<�            ����    @   �            D\�           l���0��<�    D       ����    @   \�            h��           ����0��<�    h       ����    @   ��            ��           �(�0��<�    �       ����    @   �            �X�           h�p�    �        ����    @   X�            ���           ����<�    �       ����    @   ��            ���           ���    �        ����    @   ��            4�           D�L�            ����    @   4�            H|�           ����    H        ����    @   |�            x��           ����    x        ����    @   ��            ��           �$�    �        ����    @   �            �T�           d�l�    �        ����    @   T�            ���           ����    �        ����    @   ��            0��           �� ��    0       ����    @   ��            L0�           @�L��    L       ����    @   0�            h|�           �����    h       ����    @   |�            ���           �����    �       ����    @   ��            ��           $�0��    �       ����    @   �            �`�           p�|��    �       ����    @   `�            ���           �����    �       ����    @   ��            ���           ���    �       ����    @   ��            D�           T�`�<�           ����    @   D�            8��           �����    8       ����    @   ��            X��           �����    X       ����    @   ��            x(�           8�D��    x       ����    @   (�            �t�           ������<�    �       ����    @   t�            ���           ����    �        ����    @   ��            ��           �$�    �        ����    @   �             T�           d�t��<�            ����    @   T�            8��           ����<�    8       ����    @   ��            X��            ��<�    X       ����    @   ��            p<�           L�T�    p        ����    @   <�            ���           ����    �        ����    @   ��            ���           ���������<�    �       ����    @   ��            L��            �8�           H�\����<�    �       ����    @   8�            ��           ����\����<�           ����    @   ��            ����            D��           ��H�    D       ����    @   ��            dD�           T�d��<�    d       ����    @   D�            ���           �����<�    �       ����    @   ��            ���           ��� ��<�    �       ����    @   ��            �8�           H�X��<�    �       ����    @   8�            ���           �����<�    �       ����    @   ��             ��           �������<�            ����    @   ��            $,�           <�P����<�    $       ����    @   ,�            H��           �������<�    H       ����    @   ��            l��           �������<�    l       ����    @   ��            �(�           8�L����<�    �       ����    @   (�            �|�           �����<�    �       ����    @   |�            ���           ����    �        ����    @   ��            ��           $�4��<�    �       ����    @   �            d�           t����<�           ����    @   d�            (��           �������<�    (       ����    @   ��            � ��            D�           ,�@����<�    D       ����    @   �            dp�           �������<�    d       ����    @   p�            ���           ���������<�    �       ����    @   ��            ��(�            �0�           @�L�<�    �       ����    @   0�            �|�           ����<�    �       ����    @   |�            ���           ������<�    �       ����    @   ��            ��           (�4�<�    �       ����    @   �            d�           t���4�<�           ����    @   d�            4��           ������4�<�    4       ����    @   ��            X             ( 4�<�    X       ����    @                xX            h p     x        ����    @   X             ��            � �     �        ����    @   �             ��            �      �        ����    @   �             �0           @P��<�    �       ����    @   0            �           ��<�           ����    @   �            ,�           ��    ,        ����    @   �            `           $,    `        ����    @               �\           lx<�    �       ����    @   \            ��           ���    �       ����    @   �            ��           ��    �       ����    @   �            D           T`,           ����    @   D            4�           ��`,    4       ����    @   �            X�           � ��<�    X       ����    @   �            �0           @L<�    �       ����    @   0            �|           ����,�    �       ����    @   |             �           ��             ����    @   �            ����            d&(           8D��    d&       ����    @   (� �� @: Ԓ �� d  �  ! M! �! �" �" 1# [# �# �$ �$ % �% �% �% 
& �+ �+ �+ (, X, �, �, �, J- j. �. �. ./ _/ �/ �1 !2 Q2 �2 �2 �2 3 H3 x3 �3 �3 4 84 h4 �4 �4 �5 �5  6 .6 ^6 �6 �6 �6 7 V7 �7 �7 �7 +8 [8 �8 �8 �8 19 X9 �9 %: K: {: �: �: ; H; {; �; < 8< h< �< �< = ;= h= �= �=  > (> n> �> �> �> (? [? �? �? �? @ H@ x@ �@ �@ !A qA �A �A LB xB �B �B 8C kC �C �C D ID {D �D �D E ;E kE �E �E �E +F aF �F �F �F FG �G �G �G +H [H �H �H �H 6I &J K KK {K �K �L �L �M �M &N XN �N �N O ;O kO �O �O �O (P �P CQ hQ �Q �Q $R KR {R �R �R S KS �S �S T \T �T �T �T ;U �U �U �U V VV �V �V 1W aW �W �W X gX Y HY xY �Y �Y Z ;Z �Z �Z [ \[ �[ �[ \ H\ �\ �\ �\ ] S] �] �] �] (^ q^ �^ �^ _ >_ �_ �_ �_ m` �` �` a 8a ha �a �a  b Qb {b �b �b c ;c kc �c �c �c +d [d �d 1e ae �e �e �e �f g @g �g �g <h ph �h �h �h (i Xi �i �i �i +j [j �j k Hk {k �k �k l ;l hl �l �l �l 1m am �m �m �m !n Qn �n �n �n o Ho xo �o p Xp �p �p �p q Kq �q �q �q +r kr �r �r s ;s �t �u v qv �v +w Xw qx �x �x y ;y �y �y �y 1z cz �z �z �z { K{ {{ �{ | I| {| �| �| } K} x} �} �} ~ ;~ h~ �~ �~ �~ ( X � � � �� ˀ � F� x� �� � 1� �� � Y� �� �� �� O� {� х � H� {� �� � !� Q� {� �� � � I� �� �� ؈ � A� q� �� Ӊ  � i� �� � � 3� �� �� �� � K� {� �� ۍ ,� a� �� ێ � Y� ݏ � K� x� � P� �� ȑ �� �� �� �� 0� X� �� �� � ]� �� ɔ �� 3� v� �� ە )� c� �� Ö �� L� �� ̗ �� 9� h� �� ۘ  � H� x� �� ؙ � 8� �� ۚ � ;� k� �� ț �� >� y� �� � � X� �� �� � #� S� �� �� � 9� h� �� � _� �� � 1� k� �� ء � ;� �� ܢ S� �� � 1� p� �� � � �� ȥ � >� h� �� � ,� |� �� � � K� �� � z�  � P� �� Ϊ �� (� X� �� �� � � K� {� �� � &� X� �� �� � � H� x� �� � � 8� v� �� د � ;� k� �� ˰ �� +� X� �� �� � � K� {� �� ۲ /� X� �� ȳ � 8� v� �� � � H� �� �� � @� v� �� ض � 8� k� �� ˷ �� +� [� �� �� � � K� {� �� � � K� �� Ժ � (� X� �� �� � � H� x� �� ؼ � 8� h� �� Ƚ �� 3� y� �� ؾ � ;� k� �� ˿ �� +� [� �� �� �� � H� x� �� �� � C� h� �� �� �� +� [� �� �� �� +� [� �� �� �� #� ^� �� �� �� � K� {� �� � H� {� �� �� � Y� �� �� �� ;� �� �� � P� �� �� � H� �� �� �� � K� �� �� I� {� �� �� � 8� ~� �� �� � K� �� �� � 8� h� �� �� � _� �� �� +� X� �� �� �� � K� {� �� �� =� �� �� � ;� k� �� �� �� +� [� �� �� �� !� K� x� �� 8� �� � ;� s� �� �� �� >� ~� �� � K� {� �� � >� s� �� �� � H� x� �� �� � I� �� �� �� <� h� �� �� �� (� �� ��  � (� i� �� �� � C� s� �� �� !� �� �� �� � a� �� &� [� �� �� +� `� �� �� �� )� `� �� �� �� � }� �� &� X� �� �� �� � S� �� �� �� � ;� h� �� �� �� +� [� �� �� �� (� X� �� �� �� � H� x� �� �� (� f� �� �� � V� �� �� � O� �� �� � ;� k� �� �� �� +� X� �� �� � @� s� �� ?� �� �� �� � ;� s� �� �� �� +� a� �� �� �� +� [� �� )� c� �� �� � .� Q� l�                     "�   �                       ����0     8    C    N    Y "�                           �����     �    �    �    � "�   L                       �����     �    �    �    !   	!   !����4!"�   �                       ����p!"�   �                       "�                           �����!    �!   �!   �!   �!   �!   �!   �!   �!   "	   "
   "   ""   -"   8"   C"   N"   Y"   d"   o"   w"   �"   �"   �"   �"�����"    �""�   �                       ����#    #"�   �                                 @   Lh    h�    ����       ��     ��    ����       h�����P#"�   �                       ����y#"�   �                       "�#                           �����#    �#   �#   �#   �#   �#   �#   �#   �#    $	   $   $   $   $   $   $   $   $   $   $   $   &$   .$   6$   A$   I$   Q$   Y$   d$   o$   z$   �$   �$    �$!   �$�����$    �$   �$"�                          ����%    
%   %"�   T                       "�   �                       ����;%    C%    N%   V%    ^%   f%    n%   v%    ~%   �%    �%�����%    �%"�                          �����%"�   @                       ����&"�   l                       "�   �                       ����%&    0&   ;&   F&   Q&   \&   g&   r&   }&   �&   �&
   �&   �&   �&   �&   �&   �&   �&   �&   �&   �&   	'   '   '   *'   2'   ='   H'   S'   ^'   i'   t'   '    �'   �'"   �'   �'$   �'   �'&   �'   �'(   �'   �'*   �'   (,   (   (.   $(   /(0   :(   E(2   P(   [(4   f(   q(6   |(   �(8   �(   �(   �(;   �(   �(=   �(>   �(=   �(@    )=   )B   )=   !)D   ,)=   7)F   B)=   M)H   X)=   c)J   n)=   y)L   �)=   �)N   �)=   �)P   �)=   �)R   �)=   �)T   �)=   �)V   �)=   �)X   *=   *Z   *=   )*\   4*=   ?*^   J*=   U*`   `*=   k*b   v*=   �*d   �*=   �*f   �*=   �*h   �*=   �*j   �*=   �*=   �(m   �(m   �*o   �*m   �*q   +m   +s   +m   #+u   .+m   9+w   D+m   O+y   W+z   b+y   m+y   x+}   �+@           ګ @           k� ����    ����                  "�   �                              �              ������+"�   @                       ���� ,"�   l                            �     �����P,"�   �                          � h    ��    ����    (   ��     ��    ����    (   � �����,"�                          �����,"�   H                       �����,"�   t                       ����-    )-   1-"�   �                       "�#                            ����e-    m-   u-   }-   �-   �-   �-   �-   �-   �-	   �-   �-   �-   �-   �-   �-   �-   �-   �-   �-   �-   �-   �-   �-    .   .   .   .   #.   ..   9.   D.   O.    W.!   b.�����.    �.   �."�   !                       �����."�   T!                       "�
   �!                       �����.�����.   �.   �.   �.   /   /   /   /   &/����L/    W/"�   �!                       ����}/�����/   �/"�   ("                       "�*   �"                       �����/    �/    �/    �/    �/    �/   �/    0   0   0	   '0	   I0   T0   _0   j0   u0	   �0	   �0   �0   �0   �0   �0   �0   �0   �0   �0   1   !1   ,1   41   S1   ^1   i1    t1!   1"   �1#   �1   �1%   �1%   �1'   �1'   �1����2"�   �#                       ����@2"�   $                       ����p2"�   0$                       �����2"�   \$                       �����2"�   �$                       ���� 3"�   �$                       ����@3"�   �$                       ����p3"�   %                            �     t%�����3"�   H%                          �% h    P�    ����    (   ������3"�   �%                       ���� 4"�   �%                       ����04"�   �%                       ����`4"�   $&                       �����4"�   P&                       �����4    �4"�   |&                       "�   �&                       ���� 5    5����5   !5   ,5   N5   p5   {5�����5"�   '                       �����5    �5"�   @'                       ���� 6"�   t'                       ����P6"�   �'                       �����6"�   �'                       �����6"�   �'                       �����6"�   $(                       ����7"�   P(                       ����@7    H7"�   |(                       �����7"�   �(                       �����7    �7   �7"�   �(                       �����7"�   )                       ���� 8"�   D)                       ����P8"�   p)                       �����8    �8   �8"�   �)                       �����8"�   �)                       �����8"�   *                       ���� 9"�   0*                       ����P9"�   \*                       "�   �*                       �����9    �9   �9   �9   �9"�   �*                       �����9    �9   �9   �9   	:   :����@:"�   (+                       ����p:"�   T+                       �����:"�   �+                       �����:"�   �+                       ����;"�   �+                       ����@;"�   ,                       ����p;"�   0,                       �����;�����;�����;"�   \,                       �����;    �;����<"�   �,                       ����0<"�   �,                       ����`<"�    -                       �����<�����<"�   ,-                       �����<�����<"�   `-                       ���� ="�   �-                       ����0="�   �-                       ����`="�   �-                       �����="�   .                       �����="�   D.                       �����=�����="�   p.                       ���� >"�   �.                       ����P>    [>   c>"�   �.                       �����>"�   /                       �����>"�   8/                       �����>"�   d/                       ���� ?"�   �/                       ����P?"�   �/                       �����?"�   �/                       �����?"�   0                       �����?"�   @0                       ����@"�   l0                       ����@@"�   �0                       ����p@"�   �0                       �����@"�   �0                       �����@"�   1                       ���� A    A   A"�   H1                       ����PA    [A   fA"�   �1                       �����A    �A   �A   �A"�   �1                       �����A"�   2                       ���� B    +B����6B����AB"�   02                       ����pB"�   t2                       �����B�����B   �B   �B"�   �2                       �����B"�   �2                       ����0C"�   3                       ����`C"�   <3                       �����C"�   h3                       �����C"�   �3                       ���� D"�   �3                       ����0D"�   �3                       ����pD"�   4                       �����D"�   D4                       �����D"�   p4                       ���� E"�   �4                       ����0E"�   �4                       ����`E"�   �4                       �����E"�    5                       �����E"�   L5                       �����E"�   x5                       ���� F"�   �5                       ����PF"�   �5                       �����F"�   �5                       �����F    �F"�   (6                       �����F"�   \6                       ����0G    8G"�   �6                       ����pG    {G   �G   �G"�   �6                       �����G"�    7                       �����G"�   ,7                       ���� H"�   X7                       ����PH"�   �7                       �����H"�   �7                       �����H    �H"�   �7                       �����H"�   8                       ���� I����+I"�   <8                       "�   �8                       ����`I    hI   sI   ~I   �I   �I   �I   �I   �I   �I	   �I
   �I   
J   J"�   (9                       ����PJ    XJ   cJ   nJ   yJ   �J   �J   �J   �J   �J	   �J
   �J   �J   K����@K"�   �9                       ����pK"�   �9                       �����K"�   �9                       "�   @:                       �����K    �K   �K   �K   �K   L   L    L   .L   FL	   ^L
   lL   zL   �L�����L"�   �:                       "�    ;                       �����L    �L   M   M   M   $M   2M   @M   NM   fM	   ~M
   �M   �M   �M�����M"�   p;                       ����N    N"�   �;                       ����PN"�   �;                       �����N"�   �;                       �����N    �N"�   (<                       �����N    �N"�   \<                       ����0O"�   �<                       ����`O"�   �<                       �����O"�   �<                       �����O"�   =                       �����O"�   @=                       ���� P"�   l=                       "�
   �=                       ����PP    XP   cP   nP   yP   �P   �P   �P   �P   �P"�	   0>                       �����P    �P   �P   �P   	Q   Q   Q   *Q   5Q����`Q"�   x>                       �����Q�����Q"�   �>                       �����Q    �Q   �Q"�   �>                       ���� R    R   R"�   ?                       ����@R"�   P?                       ����pR"�   |?                       �����R"�   �?                       �����R    �R"�   �?                       ���� S����S"�   @                       ����@S"�   <@                       ����pS����xS   �S"�   h@                       �����S"�   �@                       �����S    �S   �S   �S"�   �@                       ����0T    8T   CT   NT"�   A                       �����T"�   XA                       �����T"�   �A                       �����T    �T"�   �A                       ���� U    (U   0U"�   �A                       ����yU    `U"�    B                       �����U"�   TB                       �����U"�   �B                       ����V"�   �B                       ����@V    KV"�   �B                       "�   0C                       �����V�����V�����V�����V�����V�����V"�   XC                       ���� W"�   �C                       ����PW"�   �C                       �����W"�   �C                       �����W"�   D                       �����W    �W   �W   �W"�   4D                       "�   �D                       ����0X    ;X    CX   NX   YX"�   �D                       �����X    �X   �X   �X   �X   �X   �X   �X   �X    �X    Y����@Y"�   @E                       ����pY"�   lE                       �����Y"�   �E                       �����Y"�   �E                       ���� Z"�   �E                       ����0Z"�   F                       ����`Z    kZ   vZ   �Z"�   HF                       �����Z�����Z�����Z"�   �F                       �����Z    �Z"�   �F                       ����0[    ;[   F[   Q["�   �F                       �����["�   @G                       �����["�   lG                       �����[    �["�   �G                       ����@\"�   �G                       ����p\    x\"�   �G                       �����\    �\"�   ,H                       �����\"�   `H                       ����]"�   �H                       ����@]    K]"�   �H                       �����]    �]"�   �H                       �����]"�    I                       �����]"�   LI                       ���� ^"�   xI                       ����P^    X^   c^"�   �I                       �����^    �^"�   �I                       �����^    �^"�   J                       �����^    �^"�   HJ                       ���� _    (_   3_"�   |J                       ����`_    h_   s_   ~_"�   �J                       �����_    �_"�   �J                       �����_"�   0K                       "�   �K                       ���� `����+`   6`   A`����L`   b`�����`    �`"�   �K                       �����`"�   �K                       ���� a"�   L                       ����0a"�   <L                       ����`a"�   hL                       �����a"�   �L                       �����a    �a   �a   �a"�   �L                       ���� b    b   b   b"�   M                       ����@b"�   HM                       ����pb"�   tM                       �����b"�   �M                       �����b"�   �M                       ���� c"�   �M                       ����0c"�   $N                       ����`c"�   PN                       �����c"�   |N                       �����c"�   �N                       �����c"�   �N                       ���� d"�    O                       ����Pd"�   ,O                       "�   |O                       �����d�����d�����d   �d�����d   �d�����d   �d�����d   �d�����d
   �d���� e"�   �O                       ����Pe"�   P                       �����e"�   4P                       �����e"�   `P                       �����e"�   �P                       "�
   �P                       ����f    f   #f   .f   9f   Df   Of   Zf   ef   sf"�
   PQ                       �����f    �f   �f   �f   �f   �f   �f   �f   �f   g����0g    8g"�   �Q                       ����`g    kg   vg   �g"�   �Q                       �����g    �g   �g   �g"�   R                       "�   �R                       ���� h    h   h   h   &h   1h����`h    hh"�   �R                       �����h        "�   �R                       �����h"�   S                       �����h        "�   DS                       ���� i"�   xS                       ����Pi"�   �S                       �����i"�   �S                       �����i�����i�����i�����i"�   �S                       �����i"�   @T                       ���� j"�   lT                       ����Pj"�   �T                       "�
   �T                       �����j    �j   �j   �j   �j   �j   �j   �j   �j   �j����k"�   8U                       ����@k"�   dU                       ����pk"�   �U                       �����k"�   �U                       �����k"�   �U                       ���� l"�   V                       ����0l"�   @V                       ����`l"�   lV                       �����l"�   �V                       �����l"�   �V                       �����l"�   �V                       ���� m"�   W                       ����Pm"�   HW                       �����m"�   tW                       �����m"�   �W                       �����m"�   �W                       ����n"�   �W                       ����@n"�   $X                       ����pn"�   PX                       �����n"�   |X                       �����n"�   �X                       ���� o"�   �X                       ����0o����8o����@o"�    Y                       ����po"�   <Y                       "�   �Y                       �����o    �o   �o   �o   �o   �o����p"�   �Y                       ����Pp"�   �Y                       �����p"�   Z                       �����p"�   @Z                       �����p"�   lZ                       ����q"�   �Z                       ����@q"�   �Z                       �����q"�   �Z                       �����q"�   [                       �����q"�   H[                       ���� r"�   t[                       ����`r"�   �[                       "�   �[                       ����    ����    ����    ����    ����    ����    ����    �����r����           ����    ����    ����    �����r����    ����    �����r"�   p\                       ���� s"�   �\                       ����0s"�   �\                       "�   ]                       ����ps    {s   �s   �s   �s   �s   �s   �s   �s   �s	   �s
   t   t    t   .t   <t   Jt   Xt   ft   tt   �t   �t"�   �]                       �����t    �t   �t   �t   �t    u   u   u   *u   8u	   Fu
   Tu   bu   pu   ~u   �u   �u   �u   �u   �u   �u   �u����v"�   �^                       ����Pv����[v����fv"�   �^                       "�   (_                       �����v    �v   �v   �v   �v   �v   �v���� w"�   `_                       ����Pw"�   �_                       "�   �_                       �����w�����w�����w�����w�����w�����w�����w�����w�����w�����w�����w����x����x����!x   ,x����7x����Ex����Px����[x����fx�����x    �x"�   |`                       �����x"�   �`                       ���� y"�   �`                       ����0y"�   a                       "�   Xa                       ����`y    ky   vy    vy   �y�����y    �y"�   �a                       �����y    �y"�   �a                       ����z    z   #z"�   �a                       ����Pz    Xz"�   $b                       �����z"�   Xb                       �����z"�   �b                       �����z"�   �b                       ����{"�   �b                       ����@{"�   c                       ����p{"�   4c                       �����{"�   `c                       "�   �c                       �����{    �{   �{   �{   �{���� |    (|   3|   >|"�   �c                       ����p|"�   d                       �����|"�   Hd                       �����|"�   td                       ���� }"�   �d                       ����0}����8}   @}"�   �d                       ����p}"�   e                       �����}"�   4e                       �����}"�   `e                       ���� ~"�   �e                       ����0~"�   �e                       ����`~"�   �e                       �����~"�   f                       �����~"�   <f                       �����~"�   hf                       ���� "�   �f                       ����P"�   �f                       �����"�   �f                       �����    �   �"�   g                       ���� �"�   Tg                       "�
   �g                       ����0�    ;�   F�   Q�   \�   g�   r�   }�   ��   ��������"�   �g                       ������    ��"�    h                       ����0�    8�"�   Th                       ����p�"�   �h                       ������"�   �h                       ����Ё    ہ   �   �"�   �h                       ���� �"�   $i                       "�   ti                       ����P�    X�   f�   t�   ��   ��   ��"�   �i                       ����Ђ    ؂   �   �   �   �����@�����H�"�    j                       ������"�   4j                       ������"�   `j                       "�   �j                       ������    �   �   �   �   �   +�   9�   G�   U�	   c�
   q�   �"�   <k                       ������    ��   Ä   ф   ߄   �   ��   	�   �   %�	   3�
   A�����p�"�   �k                       ����������������ƅ"�   �k                       ���� �"�   l                       ����@�"�   0l                       ����p�"�   \l                       ������    ��"�   �l                       ������"�   �l                       �����"�   �l                       ����@�"�   m                       ����p�"�   @m                       ������"�   lm                       ����Ї"�   �m                       ���� �"�   �m                       ����0�    ;�"�   �m                       ����p�    x�"�   $n                       ������    ��"�   Xn                       ����Ј"�   �n                       ���� �"�   �n                       ����0�"�   �n                       ����`�"�   o                       ������"�   <o                       ������    ȉ"�   ho                       "�   �o                       ���� ������������������   ����������@�    H�   S�   ^�"�   �o                       ������    ��"�   4p                       "�   �p                       ������    ��    	�    �    �"�   �p                       ����0�    ;�    I�    T�    b�   m�    x�    ��   ��    ��    ��
   ��    ��    ΋   ً���� �    (�"�   Pq                       ����p�    x�    ��        "�   �q                       ������    ��"�   �q                       ������    �"�   �q                       �����"�   0r                       ����@�"�   \r                       ����p�"�   �r                       ������"�   �r                       ����Ѝ"�   �r                       ���� ���������������$�"�   s                       ����P�"�   Ps                       ������������   ��"�   |s                       ����Ў"�   �s                       �����"�   �s                       ����@�    K�"�   t                       "�   ht                       ����������������������������������Ǐ����ҏ�����"�   �t                       ����@�"�   �t                       ����p�"�   �t                       "�	   Hu                       ������    ��   ��   ��   ̐   א   �   �   ��"�   �u                       ���� �    (�����0�   8�����@�   H�"�   v                       ����p�    x�������   ��������   ��������"�   8v                       �����"�   dv                       "�
   �v                       ���� �    +�   6�   A�   L�   W�   b�   m�   x�   ��������"�   w                       ������"�   0w                       ���� �    (�"�   \w                       ����P�"�   �w                       ������"�   �w                       ������"�   �w                       ������"�   x                       "�   dx                       �����    �   &�   1�   <�   G�   R�������"�   �x                       ������"�   �x                       �����"�   �x                       ���� �    (�"�    y                       ����P�����[�����f�����n�"�   Ty                       ������"�   �y                       ����Е"�   �y                       ���� �    �   �   �"�   �y                       ����P�    X�"�   4z                       ������"�   hz                       ������    ��"�   �z                       ������    �   �"�   �z                       ���� �    (�   3�   >�"�   {                       ����p�    x�"�   H{                       ������    ��   ��   ��"�   |{                       �����"�   �{                       ���� �"�   �{                       ����`�"�   |                       ������������"�   D|                       ����И"�   x|                       ���� �    �   �   �"�   �|                       ����@�"�   �|                       ����p�"�   }                       ������    ��"�   @}                       ����Й"�   t}                       ���� �    �"�   �}                       ����0�"�   �}                       "�   $~                       ����`�����h�   p�   x�   ��   ��������    ˚   Ӛ"�   T~                       ���� �"�   �~                       ����0�"�   �~                       ����`�"�   �~                       ������"�                          ������"�   @                       �����"�   l                       ���� �    +�����3�"�   �                       ����`�"�   �                       ������"�    �                       ����М    ۜ   �"�   ,�                       �����"�   h�                       ����@�    H�   P�"�   ��                       ������"�   Ѐ                       ������"�   ��                       ������"�   (�                       �����    �"�   T�                       ����@�    H�"�   ��                       ����p�    x�   ��"�   ��                       ������"�   ��                       ������"�   $�                       �����    �   #�   .�"�   P�                       ����`�"�   ��                       ������    ��   ��"�   ��                       ������    �   ��"�   ��                       ����0�    ;�    F�   Q�"�   8�                       ������    ��������"�   |�                       ����Р    ۠    �"�   ��                       �����    �   &�"�   �                       ����`�"�   0�                       ������"�   \�                       ����С"�   ��                       ���� �"�   ��                       ����0�"�   ��                       "�   0�                       ����`�    h�   s�   ~�   ��������    ��   Ƣ   Ѣ"�   X�                       "�   ��                       ���� �    �   �   !�   ,�   7�   E�"�   �                       ������    ��   ��   ��   �������"�   D�                       �����    �   &�"�   p�                       ����`�    h�"�   ��                       ������    ��"�   ��                       ����Ф    ؤ"�   �                       ���� �    �"�   H�                       "�   ��                       ����0�����8�   @�   K�   S�   [�����c�����k�   s�   ~�	   ��	   ��������"�    �                       �����    ��"�   ,�                       ���� �    (�   3�"�   `�                       ����`�"�   ��                       ������"�   Ȉ                       ����Ц    ئ"�   �                       ���� �    �    �    !�"�   (�                       ����P�    [�   f�   q�"�   l�                       ������    ��"�   ��                       �����"�   �                       �����"�   �                       ����@�"�   <�                       "�   ��                       ����p�    x�    ��   ��    ��   ������Ш    ب   �   �"�   ��                       "�	   $�                       ���� �    (�   3�   >�   F�   N�   Y�   d�   o�"�	   ��                       ������    ��   ��   ��   é   Ω   ٩   �   �����0�    8�   @�   H�"�   ؋                       ����p�    x�   ��"�   �                       ������������   ê"�   X�                       �����"�   ��                       ���� �"�   ��                       ����P�"�   �                       ������"�   �                       ������"�   D�                       �����"�   p�                       �����"�   ��                       ����@�"�   ȍ                       ����p�"�   �                       ������"�    �                       �����"�   L�                       �����    �"�   x�                       ����P�"�   ��                       ������"�   ؎                       ������"�   �                       �����    �"�   0�                       �����"�   d�                       ����@�"�   ��                       ����p�"�   ��                       ������"�   �                       ����Ю    خ"�   �                       ���� �    �"�   H�                       ����0�"�   |�                       ����`�    h�"�   ��                       ������"�   ܐ                       ����Я"�   �                       ���� �"�   4�                       ����0�"�   `�                       ����`�"�   ��                       ������"�   ��                       ������"�   �                       �����"�   �                       ���� �"�   <�                       ����P�"�   h�                       ������"�   ��                       ������"�   ��                       �����"�   �                       �����"�   �                       ����@�"�   D�                       ����p�"�   p�                       ������"�   ��                       ����в"�   ȓ                       ���� �    �   �   !�"�   ��                       ����P�"�   8�                       ������    ��"�   d�                       ������"�   ��                       �����    ��"�   Ĕ                       ����0�"�   ��                       ����`�    k�"�   $�                       ������"�   X�                       ����д    ش"�   ��                       �����"�   ��                       ����@�"�   �                       ����p�    x�"�   �                       ������"�   D�                       �����    �   �   �"�   p�                       ����0�    8�"�   ��                       ����`�    k�"�   �                       ������"�   �                       ����ж"�   H�                       ���� �"�   t�                       ����0�"�   ��                       ����`�"�   ̗                       ������"�   ��                       ������"�   $�                       �����"�   P�                       ���� �"�   |�                       ����P�"�   ��                       ������"�   Ԙ                       ������"�    �                       �����"�   ,�                       �����"�   X�                       ����@�"�   ��                       ����p�"�   ��                       ������"�   ܙ                       ����й    ع   �"�   �                       �����"�   D�                       ����@�"�   p�                       ����p�    x�   ��"�   ��                       ������    ��   ƺ"�   ؚ                       �����"�   �                       ���� �"�   @�                       ����P�"�   l�                       ������"�   ��                       ������"�   ě                       �����"�   �                       �����"�   �                       ����@�"�   H�                       ����p�"�   t�                       ������"�   ��                       ����м"�   ̜                       ���� �"�   ��                       ����0�"�   $�                       ����`�"�   P�                       ������"�   |�                       ������"�   ��                       �����"�   ԝ                       ���� �    (�"�    �                       ����P�    X�   c�   n�"�   4�                       ������"�   x�                       ����о"�   ��                       ���� �"�   О                       ����0�"�   ��                       ����`�"�   (�                       ������"�   T�                       ������"�   ��                       �����"�   ��                       ���� �"�   ؟                       ����P�"�   �                       ������"�   0�                       ������"�   \�                       ������"�   ��                       �����"�   ��                       ����@�"�   �                       ����p�"�   �                       ������"�   8�                       ������"�   d�                       ���� �"�   ��                       ����0�    8�"�   ��                       ����`�"�   �                       ������"�   �                       ������"�   H�                       ������"�   t�                       ���� �"�   ��                       ����P�"�   ̢                       ������"�   ��                       ������    ��   ��"�   $�                       ������"�   `�                       ���� �"�   ��                       ����P�"�   ��                       ������"�   �                       ������"�   �                       ������"�   <�                       �����    �"�   h�                       ����@�    H�   S�"�   ��                       ������"�   ؤ                       ������"�   �                       ������"�   0�                       �����"�   \�                       ����@�"�   ��                       ����p�"�   ��                       ������    ��   ��"�   �                       ������    �   �"�   �                       ����@�"�   X�                       ����p�"�   ��                       ������    ��"�   ��                       ������    ��"�   �                       �����"�   �                       ����@�"�   D�                       ������"�   p�                       ������"�   ��                       ������"�   ȧ                       �����    �   #�"�   ��                       ����`�    h�   s�"�   0�                       ������"�   l�                       ������    ��   ��"�   ��                       ����0�    8�   @�   H�"�   Ԩ                       ������    ��   ��   ��"�   �                       ������"�   \�                       ���� �    �"�   ��                       ����@�"�   ��                       ����p�    x�"�   �                       ������"�   �                       ������"�   H�                       �����"�   t�                       ����@�"�   ��                       ����p�    x�   ��   ��"�   ̪                       ������������"�   �                       "�   h�                       ���� ������   ������   #�����+�����3�����>�����p�"�   ��                       ������"�   ԫ                       ������"�    �                       ���� �"�   ,�                       ����0�"�   X�                       ����`�    k�����v�"�   ��                       ������"�   ��                       ������    ��"�   �                       �����"�    �                       ����@�"�   L�                       ����p�    {�"�   x�                       ������    ��   ��"�   ��                       ���� �"�   �                       ����0�"�   �                       ����`�"�   @�                       ������"�   l�                       ������"�   ��                       ������    ��"�   Į                       "�   �                       ���� �    (�   3�   >�   I�   T�������"�   L�                       "�   ��                       ������    ��   ��   ��   ��   ��   ������ �"�   ԯ                       ����P�"�    �                       ������"�   ,�                       ������"�   X�                       ������    ��"�   ��                       �����"�   ��                       ����@�"�   �                       ����p�"�   �                       ������"�   <�                       ������"�   h�                       "�   ��                       ���� �    �   �   !�   /�"�   �                       ����`�    h�   s�   ��   ��������"�   ,�                       ������    ��"�   X�                       ����0�"�   ��                       ����`�"�   ��                       ������"�   �                       ������"�   �                       ������"�   <�                       ���� �"�   h�                       ����P�"�   ��                       ������"�   ��                       ������"�   �                       ������"�   �                       �����"�   D�                       ����@�"�   p�                       ����p�"�   ��                       ������"�   ȴ                       "�   �                       ������    ��   ��   ��   ��   �   �   *�"�	   |�                       ����`�    h�   s�   ~�   ��   ��   ��   ��   ������ �"�   ĵ                       ����0�"�   �                       ����`�    h�"�   �                       ������    ��"�   P�                       ������"�   ��                       ������"�   ��                       ���� �    (�   3�"�   ܶ                       ����`�    h�   s�"�   �                       ������    ��"�   T�                       "�   ��                       ��������������������������������������������@�"�   �                       ����p�"�   �                       ������    ��   ��   ��"�   <�                       ������    ��"�   ��                       ���� �    (�   3�"�   ��                       ����`�    h�"�   �                       ������    ��"�   $�                       ������    ��"�   X�                       ���� �"�   ��                       ����@�"�   ��                       ����p�"�   �                       ������"�   �                       ������"�   <�                       ���� �"�   h�                       ����0�"�   ��                       ����p�"�   ��                       ������������"�   �                       ������    ��"�    �                       �����    �   &�   1�"�   T�                       ����`�"�   ��                       ������"�   Ļ                       ������"�   �                       ������"�   �                       ���� �"�   H�                       "�   ��                       ����P�    X�   c�   k�   s�   {�   ��������"�   м                       ������    ��"�   ��                       ���� �"�   0�                       ����P�"�   \�                       ������"�   ��                       ������"�   ��                       ������    ��   �"�   �                       ����0�    8�"�   �                       ����`�    h�"�   P�                       ������    ��"�   ��                       ������������"�   ��                       ���� �    �"�   �                       "�   D�                       ����P�    X�����c�   k�����s�   {�������������"�   |�                       ������"�   ��                       �����"�   Կ                       ����@�����K�   V�"�    �                       ������������   ��"�   <�                       "�   ��                       ������    ��   ��   ��   �   �   �   �����P�"�   ��                       ������    ��"�   �                       "�   `�                       ������    ��   ��   ��   ������ �"�   ��                       ����P�����X�"�   ��                       ������������"�   ��                       ������"�   �                       ������"�   H�                       �����"�   t�                       ����P�    X�"�   ��                       ������"�   ��                       ������    ��"�    �                       ������"�   4�                       �����"�   `�                       "�   ��                       ����@�    H�   S�   a�   o�"�   ��                       ������    ��   ��   ��   ��   �������    �"�   ,�                       ����P�"�   `�                       ������"�   ��                       ������"�   ��                       ������"�   ��                       �����"�   �                       ����@�    H�"�   <�                       ����p�    x�"�   p�                       ������"�   ��                       ������"�   ��                       ���� �"�   ��                       ����0�"�   (�                       ����`�"�   T�                       ������"�   ��                       ������"�   ��                       ������"�   ��                       ���� �"�   �                       ����P�"�   0�                       ������"�   \�                       ������"�   ��                       ������    ��"�   ��                       ���� �"�   ��                       ����P�"�   �                       ������"�   @�                       ������    ��"�   l�                       ������"�   ��                       �����"�   ��                       ����@�"�   ��                       ����p�"�   $�                       ������"�   P�                       ������    ��"�   |�                       ���� �"�   ��                       ����P�    [�"�   ��                       ������    ��"�   �                       ������    ��   ��"�   D�                       �����"�   ��                       ����@�    H�"�   ��                       ������"�   ��                       ������    ��   ��"�   �                       ���� �"�   H�                       ����0�"�   t�                       ����p�    x�"�   ��                       ������    ��"�   ��                       ������������"�   �                       ����0�"�   <�                       ����`�"�   h�                       ������"�   ��                       ������"�   ��                       ������"�   ��                       ���� �"�   �                       ����P�"�   D�                       ������    ��   ��"�   p�                       ������"�   ��                       ���� ������"�   ��                       ����0�    8�"�   �                       ����`�����h�"�   @�                       ������������"�   t�                       "�   ��                       ���� �    �    �    �    )�   4�����`�    h�����p�   x�"�   ��                       ������"�   @�                       ������"�   l�                       ���� �"�   ��                       ����0�"�   ��                       ����`�    h�"�   ��                       ������    ��"�   $�                       ������"�   X�                       ������"�   ��                       ���� �"�   ��                       ����P�"�   ��                       ������"�   �                       ������    ��"�   4�                       ������"�   h�                       ���� �"�   ��                       ����P�"�   ��                       ������"�   ��                       "�   <�                       ������    ��   ��   ��   ��   ��   ��   ��   �   �	   �����P�    X�"�   ��                       ������"�   ��                       ������    ��   ��   ��"�   ��                       ���� �"�   8�                       ����&�"�   d�                       ����I�"�   ��                           ����    ����    ������    ����    ����    ����    o�    ����    ����    ����    ͠    ����    ����    ����    �    ����    ����    ����    �    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����G�p�    ����    ����    ����    ͷ    ����    ����    ����    2�    ����    ����    ����    ��    ����    ����    ����    4�    ����    ����    ����    [�    ����    ����    ����    <�    ����    ����    ����    ��        ������    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    G�    ����    ����    ����    ��    ����    ����    ����    ,�    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    g�q�����    ����    ����N�W�@           .�����    ����                  �"�   �   ,�                   ����    ����    ����    f�    ��������    ����    ����M�Q�    ����    ����    ��������    �    ��   ��h    d&    ����       ��    ����    ����    ����    !�    ����    ����    ����    ������    ������    ����    ��������    ����    ����    ����7 ;     ����    ����    �����4�4    ����    ����    ����    �=    ����    ����    ����    Xt    ����    ����    ����    D{    ����    ����    ����    
}        A|����    ����    ����    ��    ����    ����    ����    7�    ����    ����    ����    ��    ����    ����    ����    V�    ����    ����    ����    ��    ����    ����    ����    ٠    ����    ����    ����    ��    ����    ����    ����N�j�    ����    ����    ����9�M�    ����    ����    ����    3�    ����    ����    �����6�    ����    ����    ��������    ����    ����    ����    }���         �� T! \�         b�   ��         �� \! T�         ��   L�         ��                        ��     ��     Z� f� z� �� �� �� �� �� � � "� 2� >� P� `� n� �� �� �� �� �� �� �� �� � � $� 0� H� `� j� v� �� �� �� �� �� �� �� �� D� 
� $� <� V� l� �� �� �� �� �� �� �� �  � 0� F� V� d� v� �� �� �� �� �� �� �� � � ,� B� R� .� � � �� �� �� �� ��     ��     p� |�     �UuidCreate  RPCRT4.dll  � FindClose ; CompareStringW  : CompareStringA  ELCMapStringW  DLCMapStringA  �GetSystemInfo �OutputDebugStringA  }GetModuleFileNameA  �RtlUnwind ^TerminateProcess  BGetCurrentProcess nUnhandledExceptionFilter  JSetUnhandledExceptionFilter 9IsDebuggerPresent �RaiseException  FGetCurrentThreadId  GetCommandLineA HeapFree  �GetVersionExA HeapAlloc �GetProcessHeap  qGetLastError  fGetFileType � FindFirstFileA  HeapReAlloc HeapSize  �ReadFile  � DeleteCriticalSection �GetSystemTimeAsFileTime �GetProcAddress  GetModuleHandleA  � ExitProcess � FindNextFileA VSleep GetCPInfo ,InterlockedIncrement  (InterlockedDecrement  � GetACP  �GetOEMCP  ?IsValidCodePage eTlsGetValue cTlsAlloc  fTlsSetValue dTlsFree (SetLastError  �WriteFile �GetStdHandle  $SetHandleCount  �GetStartupInfoA � FreeEnvironmentStringsA UGetEnvironmentStrings � FreeEnvironmentStringsW �WideCharToMultiByte WGetEnvironmentStringsW  HeapDestroy HeapCreate  �VirtualFree �QueryPerformanceCounter �GetTickCount  CGetCurrentProcessId QLeaveCriticalSection  � EnterCriticalSection  �VirtualAlloc  uMultiByteToWideChar 7SetStdHandle  4 CloseHandle SetFilePointer  "GetConsoleCP  3GetConsoleMode  � FlushFileBuffers  RLoadLibraryA  #InitializeCriticalSection �GetStringTypeA  �GetStringTypeW  tGetLocaleInfoA  S CreateFileA �WriteConsoleA 5GetConsoleOutputCP  �WriteConsoleW SetEndOfFile  KERNEL32.dll  *ReleaseDC GetDC USER32.dll  � EnumFontFamiliesExW GDI32.dll %GetUserNameW  ADVAPI32.dll        �YU    �          �� ��  � � �   rhinoio.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �#�#�    .?AVCommandData@@   �    .?AVBaseData@@  �    .?AVRhinoRegistrationCommand@@  �#�    .?AVbad_alloc@std@@ �    .?AVexception@std@@ �    .?AVNodeData@@  �    .?AV?$ON_SimpleArray@VON_3dPoint@@@@    �    .?AV?$ON_SimpleArray@H@@    �    .?AV?$ON_SimpleArray@N@@    �    .?AV?$ON_SimpleArray@PBVON_Mesh@@@@ �    .?AV?$ON_SimpleArray@PBVON_Curve@@@@    �    .?AVSceneLoaderData@@   �    .?AVRhinoLoaderData@@   �    .?AVlogic_error@std@@   �    .?AVlength_error@std@@  �#�    .?AVSceneSaverData@@    �    .?AVRhinoSaverData@@    �    .?AVout_of_range@std@@  �#�    .?AVRhinoSerial@@   �    .?AVSNHookClass@@   �    .?AVSHA1@@  �#�#�#�#�#�#�#�#�#�#�#�#�#�#�#�    .?AVGeSortAndSearch@@   �    .?AVNeighbor@@  �    .?AVDisjointNgonMesh@@  �#�#�#�#�    .?AVGeDialog@@  �    .?AVGeModalDialog@@ �    .?AVGeUserArea@@    �    .?AVSubDialog@@ �    .?AViCustomGui@@    �#�#�#�#�#�#�#�#�#�#�#�#�#�    .?AVC4DThread@@ �#�#�    .?AVGeToolNode2D@@  �    .?AVGeToolDynArray@@    �    .?AVGeToolDynArraySort@@    �    .?AVGeToolList2D@@  �#�#�    .?AVON_Object@@ �_Q`��A���/������W�%F�����0�                                                                                                                                                                                                                                   ����            ���������    .?AVON_UserDataHolder@@ �    .?AVON__LayerSettingsUserData@@ �    .?AVON_UserData@@   �    .?AV?$ON_SimpleArray@VON__LayerPerViewSettings@@@@  �    .?AVON__LayerExtensions@@   �    .?AV?$ON_ClassArray@VON_MaterialRef@@@@ �    .?AVON_Layer@@  �    .?AV?$ON_SimpleArray@VON_DisplayMaterialRef@@@@ �    .?AV?$ON_SimpleArray@VON_MappingChannel@@@@ �    .?AV?$ON_ClassArray@VON_MappingRef@@@@  �    .?AVON_3dmObjectAttributes@@    �3������3������3������3������3������3������3�����      �?                      �?�3������3�����      �?                              �?                              �?�3������3������3�����  �?          �?  �?              �?              �?    �3������3������3������3������3������3�����      �?                              �?                              �?  �?              �?              �?    �3������3������3������3������    .?AVON_NurbsCurve@@ �    .?AVON_Curve@@  �    .?AVON_Geometry@@   �    .?AV?$ON_SimpleArray@PAVON_Curve@@@@    �    .?AVON_CurveArray@@ �    .?AVON_MeshVertexRef@@  �    .?AVON_MeshEdgeRef@@    �    .?AVON_MeshFaceRef@@    �    .?AVON_PerObjectMeshParameters@@    �    .?AV?$ON_SimpleArray@VON_3fPoint@@@@    �    .?AV?$ON_SimpleArray@_N@@   �    .?AV?$ON_SimpleArray@VON_Color@@@@  �    .?AV?$ON_SimpleArray@UON_MeshTopologyVertex@@@@ �    .?AV?$ON_SimpleArray@UON_MeshTopologyEdge@@@@   �    .?AV?$ON_SimpleArray@UON_MeshTopologyFace@@@@   �    .?AV?$ON_SimpleArray@UON_MeshPart@@@@   �    .?AV?$ON_SimpleArray@VON_MeshFace@@@@   �    .?AV?$ON_ClassArray@VON_TextureCoordinates@@@@  �    .?AV?$ON_SimpleArray@VON_SurfaceCurvature@@@@   �    .?AV?$ON_SimpleArray@VON_2dPoint@@@@    �    .?AV?$ON_SimpleArray@VON_2fPoint@@@@    �    .?AV?$ON_SimpleArray@VON_3fVector@@@@   �    .?AVON_MeshDoubleVertices@@ �    .?AVON_Mesh@@   �    .?AVON_InstanceRef@@    �    .?AVON__IDefAlternativePathUserData@@   �    .?AV?$ON_SimpleArray@U_GUID@@@@ �    .?AV?$ON_SimpleArray@PAVON_Layer@@@@    �    .?AVON_InstanceDefinition@@ �    .?AVON__IDefLayerSettingsUserData@@ �    .?AVON_Extrusion@@  �    .?AVON_Surface@@    �    .?AVON_DisplayMeshCache@@   �    .?AV?$ON_ClassArray@VON_Extrusion_BrepForm_FaceInfo@@@@ �    .?AV?$ON_SimpleArray@UON_BrepTrimPoint@@@@  �    .?AV?$ON_ClassArray@VON_BrepVertex@@@@  �    .?AV?$ON_ClassArray@VON_BrepEdge@@@@    �    .?AV?$ON_ClassArray@VON_BrepTrim@@@@    �    .?AV?$ON_ClassArray@VON_BrepLoop@@@@    �    .?AV?$ON_ClassArray@VON_BrepFace@@@@    �    .?AV?$ON_SimpleArray@PAVON_Surface@@@@  �    .?AV?$ON_SimpleArray@VON__EDGE_ENDS@@@@ �    .?AVON_BrepVertex@@ �    .?AVON_Point@@  �    .?AVON_BrepEdge@@   �    .?AVON_CurveProxy@@ �    .?AVON_BrepTrim@@   �    .?AVON_BrepLoop@@   �    .?AVON_BrepFace@@   �    .?AVON_SurfaceProxy@@   �    .?AV?$ON_ObjectArray@VON_BrepVertex@@@@ �    .?AV?$ON_ObjectArray@VON_BrepEdge@@@@   �    .?AV?$ON_ObjectArray@VON_BrepLoop@@@@   �    .?AV?$ON_ObjectArray@VON_BrepTrim@@@@   �    .?AV?$ON_ObjectArray@VON_BrepFace@@@@   �    .?AVON_BrepVertexArray@@    �    .?AVON_BrepEdgeArray@@  �    .?AVON_BrepTrimArray@@  �    .?AVON_BrepLoopArray@@  �    .?AVON_BrepFaceArray@@  �    .?AVON_Brep@@   �    .?AVON_Light@@  �    .?AV?$ON_ClassArray@VON_UserString@@@@  �    .?AV?$ON_SimpleArray@PAVON_Bitmap@@@@   �    .?AV?$ON_ClassArray@VONX_Model_RenderLight@@@@  �    .?AV?$ON_ClassArray@VONX_Model_Object@@@@   �    .?AV?$ON_SimpleArray@PAVON_HistoryRecord@@@@    �    .?AV?$ON_ClassArray@VONX_Model_UserData@@@@ �    .?AV?$ON_SimpleArray@VON__CIndexPair@@@@    �    .?AV?$ON_ClassArray@VON_TextureMapping@@@@  �    .?AV?$ON_ClassArray@VON_Material@@@@    �    .?AV?$ON_ClassArray@VON_Linetype@@@@    �    .?AV?$ON_ClassArray@VON_Layer@@@@   �    .?AV?$ON_ClassArray@VON_Group@@@@   �    .?AV?$ON_ClassArray@VON_Font@@@@    �    .?AV?$ON_ClassArray@VON_DimStyle@@@@    �    .?AV?$ON_ClassArray@VON_HatchPattern@@@@    �    .?AV?$ON_ClassArray@VON_InstanceDefinition@@@@  �    .?AV?$ON_SimpleArray@VON_UuidIndex@@@@  �    .?AV?$ON_SimpleArray@PBVON_InstanceRef@@@@  �    .?AV?$ON_ObjectArray@VON_Linetype@@@@   �    .?AV?$ON_ObjectArray@VON_Layer@@@@  �    .?AV?$ON_ObjectArray@VON_Group@@@@  �    .?AV?$ON_ObjectArray@VON_TextureMapping@@@@ �    .?AV?$ON_ObjectArray@VON_Material@@@@   �    .?AV?$ON_ObjectArray@VON_Font@@@@   �    .?AV?$ON_ObjectArray@VON_DimStyle@@@@   �    .?AV?$ON_ObjectArray@VON_HatchPattern@@@@   �    .?AV?$ON_ObjectArray@VON_InstanceDefinition@@@@ �    .?AVONX_Model@@      �o@�    .?AVON_Texture@@    �    .?AVON_TextureMapping@@ �    .?AV?$ON_ClassArray@VON_Texture@@@@ �    .?AV?$ON_ObjectArray@VON_Texture@@@@    �    .?AVON_Material@@   ����            <	H	�    .?AVON_Viewport@@   �    .?AV?$ON_SimpleArray@VON_ClippingPlaneInfo@@@@  �    .?AV?$ON_ClassArray@VON_3dmConstructionPlane@@@@    �    .?AV?$ON_ClassArray@VON_3dmView@@@@ �    .?AV?$ON_ClassArray@VON_PlugInRef@@@@   �    .?AV?$ON_SimpleArray@VON_3dVector@@@@   �    .?AV?$ON_SimpleArray@VON_UuidPair@@@@   �    .?AVON_2dPointArray@@   �    .?AVON_3dPointArray@@   �    .?AVON_2fPointArray@@   �    .?AVON_3fPointArray@@   �    .?AVON_3fVectorArray@@  �    .?AVON_UuidList@@   �    .?AVON_UuidIndexList@@  �    .?AVON_UuidPairList@@   �    .?AVON_OBSOLETE_CCustomMeshUserData@@   �    .?AV?$ON_SimpleArray@UON_3DM_BIG_CHUNK@@@@  �    .?AVON_BinaryArchive@@  �    .?AVON_BinaryFile@@ �    .?AVON_Read3dmBufferArchive@@   �    .?AVON_TextLog@@    �    .?AVON_PolylineCurve@@  �    .?AVON_TensorProduct@@  �    .?AVON_NurbsSurface@@   �    .?AVON_SumSurface@@ �    .?AVON_SumTensor@@  �    .?AVON_RevSurface@@ �    .?AVON_RevolutionTensor@@   �    .?AVON_PolyCurve@@  �    .?AVON_UnknownUserData@@    �    .?AVON_UnknownUserDataArchive@@ �    .?AVON_DocumentUserStringList@@ �    .?AVON_UserStringList@@ �    .?AVON_TextExtra@@  �    .?AVON_DimensionExtra@@ � < >   �    .?AVON_AngularDimension2Extra@@ �    .?AVON_TextDot@@    �    .?AVON_AnnotationTextFormula@@  �    .?AVON_Annotation2@@    �    .?AVON_LinearDimension2@@   �    .?AVON_RadialDimension2@@   �    .?AVON_AngularDimension2@@  �    .?AVON_OrdinateDimension2@@ �    .?AVON_TextEntity2@@    �    .?AVON_Leader2@@    �    .?AV?$ON_SimpleArray@VON_LinetypeSegment@@@@    �    .?AVON_Linetype@@   �    .?AVON_Value@@  �    .?AV?$ON_ClassArray@VON_CurveProxyHistory@@@@   �    .?AV?$ON_SimpleArray@PAVON_Value@@@@    �    .?AV?$ON_ClassArray@VON_ObjRef@@@@  �    .?AV?$ON_ClassArray@VON_wString@@@@ �    .?AV?$ON_SimpleArray@VON_Xform@@@@  �    .?AV?$ON_ClassArray@VON_PolyEdgeHistory@@@@ �    .?AVON_BoolValue@@  �    .?AVON_IntValue@@   �    .?AVON_DoubleValue@@    �    .?AVON_PointValue@@ �    .?AVON_VectorValue@@    �    .?AVON_XformValue@@ �    .?AVON_ColorValue@@ �    .?AVON_UuidValue@@  �    .?AVON_HistoryRecord@@  �    .?AVON_StringValue@@    �    .?AVON_ObjRefValue@@    �    .?AVON_PolyEdgeHistoryValue@@   �    .?AVON_HatchExtra@@ �    .?AV?$ON_ClassArray@VON_HatchLine@@@@   �    .?AV?$ON_SimpleArray@PAVON_HatchLoop@@@@    �    .?AVON_Hatch@@  �    .?AVON_HatchPattern@@   �    .?AVON_Group@@  �    .?AV?$ON_SimpleArray@VON_OffsetSurfaceValue@@@@ �    .?AV?$ON_SimpleArray@VON_BumpFunction@@@@   �    .?AVON_OffsetSurface@@  �    .?AVON_PlaneSurface@@   �    .?AVON_ClippingPlaneSurface@@   �    .?AVON_SurfaceArray@@   �    .?AVON_PointGrid@@  �    .?AVON_PointCloud@@ �    .?AVON_AnnotationTextDot@@  �    .?AVON_AnnotationArrow@@    �    .?AVON_Annotation@@ �    .?AVON_LinearDimension@@    �    .?AVON_RadialDimension@@    �    .?AVON_AngularDimension@@   �    .?AVON_TextEntity@@ �    .?AVON_Leader@@ �    .?AVON_NurbsCage@@  �    .?AV?$ON_ClassArray@VON_Localizer@@@@   �    .?AVON_MorphControl@@   �    .?AVON_DetailView@@ �    .?AVON_LineCurve@@  �    .?AVON_CurveOnSurface@@ �    .?AVON_ArcCurve@@   �    .?AVON__OBSOLETE__CircleCurve@@ �    .?AVON_Font@@   �    .?AVON_DimStyle@@   �    .?AVON_DimStyleExtra@@  �    .?AVON_Bitmap@@ �    .?AVON_WindowsBitmap@@  �    .?AVON_WindowsBitmapEx@@    �    .?AVON_EmbeddedBitmap@@   !B c0�@�P�`�p�)�J�k���������1s2R"�R�B�r�b9��{�Z��Ӝ�����b$C4 �d�t�D�Tj�K�(�	������ō�S6r&0�v�f�V�F[�z��8�����׼��H�X�h�x@a(#8���َ��H�i�
�+��Z�J�z�jqP
3:*���˿���y�X�;���l�|�L�\",<`A�������*��h�I��~�n�^�N>2.Qp���������:�Y�x�����ʱ��-�N�o�� �0� P%@Fpg`������ڳ=���^���"�25BRwbVr�˥����n�O�,���4�$��ftGd$TDۧ������_�~��<��&�6��WfvvF4VL�m��/�ș鉊���DXeHx'h���8�(}�\�?����؛����uJTZ7jz�
��*�:.��l�Mͪ����ɍ&|ld\EL�<�,���>�]�|ߛ���ُ��n6~UNt^�.�>��    �0w,a�Q	��m��jp5�c飕d�2�����y�����җ+L�	�|�~-����d�� �jHq���A��}�����mQ���ǅӃV�l��kdz�b���e�O\�lcc=���� n;^iL�A`�rqg���<G�K���k�
����5l��B�ɻ�@����l�2u\�E���Y=ѫ�0�&: �Q�Q��aп���!#ĳV���������(�_���$���|o/LhX�a�=-f��A�vq�� Ҙ*��q���俟3Ը��x4� ��	���j-=m�ld�\c��Qkkbal�0e�N b��l{����W���ٰeP�긾�|�����bI-��|ӌeL��Xa�M�Q�:t ���0��A��Jו�=m�Ѥ����j�iC��n4F�g�и`�s-D�3_L
��|�<qP�A'�� �%�hW��o 	�f���a���^���)"�а����=�Y��.;\���l�� �������ұt9G��wҝ&���sc�;d�>jm�Zjz���	�'� 
��}D��ң�h���i]Wb��ge�q6l�knv���+ӉZz��J�go߹��ﾎC��Վ�`���~�ѡ���8R��O�g��gW����?K6�H�+�L
��J6`zA��`�U�g��n1y�iF��a��f���o%6�hR�w�G��"/&U�;��(���Z�+j�\����1�е���,��[��d�&�c윣ju
�m�	�?6�grW �J��z��+�{8���Ғ�����|!����ӆB������hn�����[&���w�owG��Z�pj��;f\��e�i�b���kaE�lx�
����T�N³9a&g��`�MGiI�wn>JjѮ�Z��f�@�;�7S���Ş��ϲG���0򽽊º�0��S���$6к���)W�T�g�#.zf��Ja�h]�+o*7������Z��-�    .?AV?$ON_SimpleArray@PAN@@  �    .?AVON_Matrix@@ �    .?AV?$ON_SimpleArray@VON_ObjRef_IRefID@@@@  �    .?AVON_MeshNgonUserData@@   �    .?AVON_BrepFaceSide@@   �    .?AV?$ON_ClassArray@VON_BrepFaceSide@@@@    �    .?AV?$ON_ClassArray@VON_BrepRegion@@@@  �    .?AVON_BrepRegion@@ �    .?AV?$ON_ObjectArray@VON_BrepFaceSide@@@@   �    .?AVON_BrepFaceSideArray@@  �    .?AV?$ON_ObjectArray@VON_BrepRegion@@@@ �    .?AVON_BrepRegionArray@@    �    .?AVON_BrepRegionTopologyUserData@@ �    .?AVON_EmbeddedFile@@   �    .?AVON_Polyline@@   (�ج       ��`�              ح          �#�#�#�    .?AVtype_info@@ N�@���D�#u�  s�              sqrt                  �?pow     asin            acos            cos             sin             atan            log             fmod         ��t������tan             log10           D�                                                                                                                                                                                                                                                                                                                                        abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     8!�  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    �#    �#�    .?AVbad_exception@std@@ ��������    ����������               ���5�h!����?      �?                                       	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                           ��   ��	   X�
   ��   ��   d�   @�   �   ��   ��   |�   D�   �   ��   ��    `�!   h�"   ��x   ��y   ��z   ���   ���   ��       ��       ���ܧ׹�fq�@      ��@�6C����?      �?exp          �"}��#  ��    �����
                                                           �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �             x   
                                                                                                                                                                                                                                                                                     ?                     
      p?  �?   _       
          �?      �C      �;      �?      �?      ���$d*d/d5d:d@dFdLdRdndsd�d�d�d�d�d�d�dee"eBeVene�e�e�e�e�e�e�ef&fFfKfefjf�f�f�f�f�f�f	gg.gBgZgng�g�g�g�g�g�g�gh2h7hQhVhvh�h�h  �����C                                                                                              �,            �,            �,            �,            �,                              �4        �p���3�,   �,8!                                                                                                                                                                                                        @�    @�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     atan2        <��������������������������   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l          ?  ?        �      ���������              �   ]   ]   ]   ]   ��   ��!   ��   ]   �\   �\   ��   ��   �\   �\    �\   �\   �\   x�   �\   p�   h�   `�   X�   P�"   L�#   H�$   D�%   <�&   0�       �D        � 0                  �i��~�@sinh         ��l��cosh         �}�!�tanh        ! ��l�A�       �            �&  ��    h�d�`�\�X�T�P��(�(�(�(�(�(�(L�H�D�@�|(<�8�4�0�,�(�$��(�(�(�(|(t(l(d(X(P(D(8( ������	         �3.   �4d�d�d�d�d�d�d�d�d��4   .      ����        ����        �p     ����    PST                                                             PDT                                                             5X5      ���5      @   �  �   ����             ��������             �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         F0�0�0�011A1f1t1�1�1�1�1�1�1&242J2c2y2�2�2�2�23"3;3E3T3o3�3�3 4484L4^4i4}4�4�4�4�4�4545L5`5x5�5�5�5�56D6v6�6�6�6�6�6&747L7d7z7�7�7�78F8W8i8r8�8�8�8�8�8�8�8�899(969L9^9g9�9�9�9�9:::Z:�:�:�:�:</<H<a<y<�<�<�<�<�<
=#=<=W=p=�=�=�=�=�=�=>)>?>"?8?    �   �23"373P3`3�3�374a4�4�4�4�4545?6v6�6�6�6�8�8�8�89&9B9]9�9�9�9�9�9:':C:Z:q:�:�:�:�:�:�:;);@;W;n;t;�;�;�;<I<�<�<�<�<�<�<�<7=j=�=>>>%>J>j>�>�>�>'?a?   0  �   0?0�0�0�1�1�1d4�4�45�5�5�678K8b8�8�89,9~9�9�9�9:+:?:�:�:�:�:�:;P;�;�;<#<j<<�<�<==/=U=f=|=	>><>�>�>�>?E?�?�?�?�?�?   @  |   0�0�0�2�2�2�2�2&3;3{3�3�3�3�3f4p4�56m6�7 88.8B8f8{8�8�8989w9�9�9�:�:2;x;�;�;4<9<Y<p<�<�<�<�<=C=]=�=>,>r>�?�?�? P  �   b0�0�02212K2i3w3�3�3�3�3414K4Y4�4�4�4j5D6�8�9:*:y:�:�:�: ;;4;K;�;�;�;�;
<7<L<h<l<p<t<�<�<�<�<�<�<==.=D=�=�=�=>:>?? `  �   S0f0|0�01K1�122�2�2�2�2�23�3 4'5>5�5�5�5�5�5�5666/696C6M6W6a6�67+7G7�7�7�7U8m8�8�8V9n9s:P;<�<�<�<�=�=H>�>?�?   p  X   !0J0p0�0�0g1�1?2�23x3�3�3�344}4�4[56�6J7b7�7e8�9�9:�:y;<`<�<8=�=:>�>??�?   �  L   0�01�1�1`2�253�3�3/4�45e5�56�8`9�97:�:�:�:g;�;�<_=e=�>}?�?�?�?�? �  �   0;1x1�1�2�23:3&4a4�455C5i5�5�5U6�6t8M9�9:-:D:]:�:�:�:�:�:�:;J;_;v;�;�;�;o<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$=(=,=0=4=8=<=@=D=H=L=P=�>�>�>   �  P   n2y2I3[3�3�3�4�4y5�5�5�566\6n6�6�6�67�7�7V8^8z8�9�9�9f;x;�;�>�>�>�>�> �  h   �1�1�1%2�2�2�2�233%3L3�3�3�3�3�344%484j4u4�;�;�;�;<8<O<f<�<�<�<�<=s=�=�=>q>�>�>�>f?{?�?�? �  �   0*0<0E0^0s0�0I1b1{1�1�1�1E2[2s2�2�2�2�2�2y3�3�34!4^4t4�45535E5X5p5�5�5�5�5�5�5�56F6W6�6�7�7�78T8�8Y9t9�9�9�9�9:P:�:�:�:�:;S;j;�;�;�;�;�;�;�;�;�; <<<(<9<T<s<   �  h   f3{3�3�3�344-4A4r4�45P5g5�5�5�516�6�7�7�7�7d8�8�8919�9�9�9':V:h:g;�;2<�<�<K=�=�=>>j>�>�?   �  p   60�0�0P1�1�2�2�2�2D3�3�3�3�3�4�455:5U5v5�5�5�5'6m6�6�7�7B9�9�9�9�9:I:f::�:�:<K<\<n<�<�<�<=3=q={=�? �  t   �0�0�0�0 1J1_1s1|1�1�1�1202L2a2�2�2�3�3�34A4R4c4y4�4�4�5�6�6�6�6�6�6�6�6�6�6�7�7�7�7�:�:;;V;c;�;�;�;<     4   &848E8L8q8X<�<�<�<==f>u>�>�>�>�>�>	?3?>?    4   �1�1�1�122v4�4�4�4�4�7�7�788f9x9�9�9�9     �   �1�1�1�3K4|4�45n5�67�7�8�8�8�8�8�8�8�8�8�8�8�8�9::::R:a:�:�:�:�:0;H;Z;�;�; <%<A<�<�<=4=M=m=�=�=�=>>I>t>�>�>�>?F?b?~?�?�? 0 �   0060K0�0�0�8$9J9X9g9�9�9�9':[:�:�:�:�:�:
;$;1;>;V;i;{;�;�;�;�;�;�;<(<D<U<h<�<�<�<�<�<�<�<==6=T=f=�=�=�=�=�=�=�= >6>R>c>v>�>�>�>�>�>�>??(?F?d?v?�?�?�?�?�?�?   @ �   000F0b0t0�0�0�0�0�0141B1O1g1y1�1�1�1�1�1�12"282T2f2x2�2�2�2�2�2333=3^3t3�3�3�3�3�344G4t4�4�4"5*545F5P5k5�5�5�5�5�56=6f6�6�67'787A7T7�7�7�788*8<8b88�8�8d9y9�9�94:B:a:q:�:�:�:�:;$;D;d;�;�;�<�<�<�<�<===H=e=�=M>�>/?Q?|?�?�?�?   P �   S0e0�0�0I1e1�1�1I2l2�2�2�2�23%3�3�3!4|4�45$5D5d5�5�5�5�56$6D6d6�6�6�6�6�6747d7�7�7�7�7$8D8t8�8�8�8$9D9d9�9�9�9�9::1:D:a:q:�:�:�:�:;A;Q;d;�;�;�;<$<A<Q<a<t<�<�<�<�<=4=_=�=�=�=�=>>4>T>>�>�>�>$?J?t?�?�?�?�?   ` �   040T0t0�0�0�01T1�1�12T2�2�2�23A3a3t3�3�3�3�34$4D4d4�4�4�4�4B5h5�5�5�5�56T6r6�6�6�6�6�6747T7t7�7�7�7 88$8D8}8�8�8�899.9C9d9~9�9�9�9�9�9:$:H:a:�:�:�:�:#;9;G;V;�;�;�;�;	<<&<T<}<�<�<�<=K=^=�=�=�=�=$>D>d>�>�>�>�>�>?1?D?�?�?�?�? p �   0$0D0d0�0�0�0�0�01!141d1�1�1�1�1�1�122Z3l3~3�3�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�5�6�67E7�7�7�7E8�8�8�89U9�9�9/:u:�:�:";U;�;�;2<e<�<�<%=U=�=�=>5>�>�>?U?�?�?�?   � �    040D0e0�0�051r1�12E2�2�2	313Y3c3�3�3�3�3454Y4�4�4�45u5�5�56-6V66�6�6&7H7�788 8p9�9�9�9;@;V;�;�;;<L<r<�<�<�<�<=e=v=�=}> � �   �1�1�1�1 22�2�2�2�342585b5h5p5�5�5�5�5,6M6S6g6n6�6�6�6�6,7M7a7/8�8�8�8�8�849�9�9�9�9�9�9�:�:�:�:;';^;w;�;<4<t<�<�<=D=�=�=�=�=>4>T>�>�>�>�?�?�?�?   � �   +0[0�01191�1�1�12$2Q2d2�2�2�2�2323Q3t3�3�3�3$4D4a4�4�4�4�45D5q5�5�5�56A6a6�6�6�6�67$7D7d7�7�7�7�7�7848T8�8�8�8l9�9�9:q:�:
;-;�;�;�;a<~<�<=.=C=�=�=>A>d>�>S?|?�?   � �   #0L0t0�01D1�1�1�1k2�23a3�3�34a4�4�4L5�5�56�6�6�6>7^7s7�7!8�8�8$9D9a9q9�9�9�9�9:4:d:�:�:�:;$;D;a;�;�;�;<0<R<�<�<�<�<=&=a=�=�=�=�=>�>�>�>�>�>�>?D?a?t?�?�?�? �   0D0d0�0�0�0�0�0'1b1�1�1�122`2�2�2�2!323T3e3s3�3�3�3�3�3�34"4D4d4�4�4�4�4�4 5545T5l5�5�5�5�5�5�5 66606m66�6�6�6�67$7D7t7�7�7�7�7�78D8d8�8�8�8�8�8$9A9T9t9�9�9�9�9::$:D:d:�:�:�:�:;$;D;d;~;�;�;�;�;�<=*=?=`=h=|=>/>K>a>�>�>�>?$?D?d?�?�?�?�?�?   � (  $0D0a0q0�0�0�0�0�0�0
11D1c1q1�1�1�1�12!212A2Q2a2t2�2�2�2�2�2�2343T3t3�3�3�3�3444g4�4�4�4�4�45575I5t5�5�5�5�5646K6_6n6~6�6�6�6�6�67747X7~7�7�7�7�7�7�78"8D8b8v8�8�8�8�8949A9Q9d9�9�9�9�9:$:D:d:�:�:�:�:;$;D;d;�;�;�;�;<$<D<l<�<�<�<=$=D=d=�=�=�=�=>$>D>d>�>�>�>�>?$?D?d?�?�?�?�? � �   0!040T0t0�0�0�0�0�01141T1v1�1�1�1�1	2*2d2�2�2�3�3�3�3�3"474�4�4�45U5�5�556�6�6%7B7W7t7�7�7�7�7818A8T8q8�8�8�8�8�89$9D9h9�9�9�9�9:4:T:t:�:�:�:�:;T;q;�;�;�;�;�;<1<O<q<�<�<�<=$=D=u=�=�=�=�=�=>$>D>Y>m>�>�>�>?d?�? � �   0D0d0�0�0�0�01$1D1t1�1�1�12$2T2t2�2�2�23A3d3�3�3�3444w4�4�4�45!5A5a5�5�5�5�56!6A6a6�6�6�6�6747T7t7�7�7�7818T8�8�8�8�8$9T9�9�9�92:Q:q:�:�:�:;1;Q;q;�;�;�;<4<d<�<�<�<�<=4=a=�=�=�=�=>>4>�>�>!?4?T?�?�?�?   �   0!0Q0t0�0�0�01$1q1�1�1�12D2d2�2�23[3�3�3�3�34D4q4�4�4�4�4�4*5D5�5�5�5
6T6t6�6R7�788*8M8�8�8�89&9O9�9�9�9�98:i:�:4;D;q;�;�;�;#<7<U<t<�<�<�<=4=T=�=�=�=�=>Q>t>�>�>�>?4?T?�?�?�?  �   0a0�0�0�0�0/1N1j1�1�1�1232a2�2�2�2�2�23F3h3~3�3�3�34#484w4�4�4�455;5P5n5*6=6u6�6�6�6�6?7h9$<=<�<�<�<�<=Z=u=H?L?P?T?�?�?�?   �   040Q0d0�0�0�0�01D1t1�1�1�1�1 3-343;3B3I3P3�3�3�3�3�3�3�3�34$4�4�4�4E5t5�5�5�5$646a6�6<7h7�7�7�78W8%9*959Z9b9�9�9�9�9!:T:�:�:;D;k;�;�;
<6<K<t<�<�<+=k=�=�= >d>�>�>�>�>?'?V?m?�?�?�? 0 �   020Q0p0�0�0�0101O1�1�1�1�12'2g2�2�2�2�2*3�3�3%4~4�45[5�5�5�5;6|6�6�6�6<7V7�7�78!8x8�8�8�849�9:t:�:�:6;H;�;�;<=<�<�<-=f=�=�=�=>/>F>t>�>�>�>?i?   @ x   0I0�0�031�1�1#2�2�2C3�3�3C4�45c5�5#6�6�6C7�7�7S8�89�9�9):s:�: ;:;`;�;�;�;$<N<�<�<=;=C=t=�=�=>Z>�>�>N?�?�?   P �   0D0�0�0�01D1�1�1�112a2�2�2�2313�3�3�3�34"4�4�4�4�5V6�6�6�6�6�6�6�6�6�6�6�7 88888888 8�8�8�89?9R9n9�9�9�9�9:4:d:�:�:�:;4;t;�;�;<1<|<�<$=D=d=�=�=�=>D>t>�>�>�>�>�>?#?7?T?d?�?�?�?�?�?�?   ` �   0"0?0K0V0t0�0�0!1A1d1�1�1 2p2�2�2�2F3t3�3�34T4n45D5�5�5�5�5`6�6�6�6�6�7�7X8�8�8�8�8�8�8�8A9�9�9�9�9
::D:d:�:(;�;	<4<d<�<�<�<-=�=>!>T>t>�>�>�>�>?4?d?�?�?   p �   00)0H0Q0�0�0�0�12E2W2s2�2�2�2 3!3=3\3x3�3�3�34 4�4�4�4�4�415?5R5p5�5�5�5�5�56'6D6�6�6�67C7�7N8z8�8�8�89D9r9�9�9:T:u:�:�:�:�:�:�:;+;K;x;�;�;�;�;�;�;�;<$<5<H<`<r<�<�>.?d?�? � �   0i0�0D1e1�1�1d2�2393�3	4�4�4�4	55,5<5Y5�5�5�5	6=6�6�6�6�6�67#7D7\7�7�7�7�7�7]9e9�9�9:':d:�:�:�:�:5;�;�;<E<�<�<%=e=�=�=5>}>�>�>?/?T?t?�?�?�?�? � �   010Q0t0�01D1N1U1\1x1�1�1242Q22�2�23$3Q3t3�3�3�34#464a4�4�4�455D5t5�5�5�56D6t6�6�6�6747Q7q7�7�7�7�7$8V8k8�89$9T9�9�9�9�;�;�;�;�<�<H>�>�>�>�>?A?Q?a?q?�?�?�?   � �   040T0w0�0�0�0�01$1A1T1�1�1�2�2*3/3�3c4v4�4#565F5�5�5�57%7b7�7�7e8�8�859u9�9:R:�:�:;U;�;�;<r<�<�<R=�=�=�=">R>�>�>(?X?l?|?�?�?   � p   0E0�0�0%1u1�12e2�23B3�3�34R4�45R5�56R6�6�657�7�7%8r8�889�95:u:�:�:5;�;�;"<e<�<=U=�=�=5>�>�>5?�?�? � �   0!0M0�0�01U1�1�1E2�2�2E3�3�354u4�4�4E5�5�5%6~6�6�607}7�7�7L8�89�9�9�9&:3:>:g:n:�:�:�:�:;; ;$;(;,;0;A;T;�;�;�;�;<!<D<d<�<�<�<�<=1=T=t=�=�=D>�> �    o7   � h   111]1�1�12e2�2�2"3R3�3�3454u4�4�425b5�5�5�5%6e6�6�6E7�7�78E8�8�8U98;[; >h>l>p>t>x>[?i?�?�?   � �   "000U0]01,1P1^1�1�1�2�2�2�2P3^3s3�3H4V4�4�45w5�5�5�5�5�5X6x6�6�6�6�6�7�7�7�7�7�7�7 8,8\8�8�8�8�8�8
9B9^9h9s9x9�9�9::K:q:�:�:�:;1;T;�;�;$<w<�<     �   Z0�0�0L2�2�23363U3h3�3�3-4�4�4f5�5]6�6#7Q7n7�7�749�9�9�:�:;D;�;�;�;<4<T<�<�<�<M=x=�=�=�=�=�=�=�=�=>>> >'>.>5><>C>J>Q>X>_>j>�>�>�>�?    T   %041@1M2R2\2�2t3y3�3�3�4	55"5F5�5�5
6\9�9:.:J:f:�:�:;�=�=�=�=�>�>�>?*?d?   �   00#0[0c0h0r0�0�0�0E1J1T1�1�1�1�1�1�1�1�1&2�2�2�2�2�2�2:3?3I3555 5Z7�7
8D8^8�8�89�9�:H;b;r;�;�;�;�;<<0<C<d<i<p<{<�<�<�<=A=�=>�>�>?Q?�?�?   0 4   0M0b0�0�2�2�2D3n3}3p4�4�4�4|5�5�5�647;�?   @    �3s5 P 8   �0�0�0R1b1�1202�2�2�2�2�2�3[4�>�>�>#?6?�?�?�?�? ` |    0D1�1�2�334�5�5�5�5�56666�6�6�6�6�6s8�8�8�8�8�8�8�8�8�8�89+9R9^9�9�9�9�9�9*;Q;b;n;w;;�;�;�;�;�;�;�;�;E<�=2>   p L   �0�0�1�12/2I2j2s2|2�2�5�6�68!8-8?8F8L8^8e8k8v8�8�8�8�8�=�=�={?�?   � l   a031@1�1�1+2C2u2�3�3)4;4s4�4�4�4�4�4�45535C5\5t5�5�5�5�6
88�8�89>9J9�9�9�9:�:�:�:�:�;�<�<L>Z>   � 0   ;0S0�0�0�02 2�2�2
313&9+959l9�9C<P<0>   � T   �3�5�5	778+8i8{8�8�8�8�8�9�9�9�9>�>�>�>�>(?/?6?=?C?R?a?t?�?�?�?�?�?�?�?�? � X   �0�0�1�12�2#323U3m3y3�3�3�3�3�34+46#6S6b6�6�6�6C7P7�7�728b8�8�8B9�9�9>:�:�:2< � @   �2�2n3�3�3`6y6E7�7�7�8�8�8r9�9:;b;<�<=;=~=�=�=N>b?   � X   0"0�0S2G3�3�3)414�4�4�4�4$5/5W5b5�5j;�;�<�<==(===V=�=�=�=>�>�>�>?V?r?�?�?   � (   %0q0:1s1�1�1s2�234B4n578*8;�; �     999�9 :�=�=     4   )0>0�1�2�2�4�4�89E9<<=<M<m<�<�<%=2=�?�?    D   1$1a3�3i4�4�4�5�56 6�7�7�7�7�7)8;8�9�9�9�:�:�:Y<k<#?6?\?x?   <   �5�5�5�5S6c6�6�67#7S7b7�7�7�7�788s8�8�8�8�8r<�=�= 0 8   �3�3M4�5�58a8i8�:!;:;_;r;�;�;C<R<�=�=�>�>Y?o?   @ L   v0�0i4~4�4�4�455&6S7b79i9~9�9<<�>�>�>�>�>�>�>�>???3?D?�?�?   P ,   90N02�2;3�7�7y:�:�:�:�;�<�<	==Y=n= ` 8   )0>0�01g233I3^3"4�4$56Y8n8::�?�?�?�?�?�?   p D   90N0f0y0�0�0�0�0�0t174M57"7�7�7�7�7�7�7
898N8�8.:�;&>=>�>!? � 4   .2@2H2Q2Z2C4T4�4�45.5=5�5�7�:�:�:�:�<�<=   � d   U0i0}0�0�0�0�0121J1q1�1�1�1�12]2�2�2�2�2�233E3U3�4�4�455�5�6�6�6�677#7L7U7^7f7U8E9>�? � `   �23�4�4�4_5d5n5�5�5�5k6p6z6�6�67�8�8�9�9�9�9	::I:[:�:�:y;�;i<{<M>`>�>�>�>�>?"?�?�?   � x   <0V0u0�0�0�0�0�122 2$2(2,20242I2[2�2�2�2�293K3�3�3�3�3)4;4y4�4�4�45+5�6�6]7b7�8�9�9C=S=g=x=c>q>�>�>?:?�?�?   � �   00G0�0�0�0+1C1�1�1�122J2�2�23P3�3�3�3-4O4q4~4�4�4�4�45P5�5�5�5$6k6K8k8�8�8�8�8�89�9:�:�:;%;|;�;�;<l<�<�< =c=s=�=>S>d>�>�>%?�? � �    0I0[0�0�0�0�0V4�5�5�5�5(6V6p6�67$7)7�7.868>8G8P8X8l8�8�8�8�8�8�8�8�9�9�9:*:3:<:D:�;�;�;�;�;�;<<<1<A<F<P<m<r<|<�<�<�<�=�=�>�>   � �   �4565I5c5v5�5�5�5�56646j6�6�6�6�6�7�788�8�8�8�8=9U99:s:�:�:�:~;�;<"<�<�<�<=1=�=�=">x>�>�>�>�>�>�>�>??"?(?C?J?P?k?r?x?�?�?�?�?�?�?�? � P   0	00e0�0�0�01a1�12P2{2�2�2+3r3�3�34(4[4�4�4�45c5�5�5d:{:"<><�>�>     L   �1�156�6�6�7�7�9�:v;};�;�;�;D<W<3=D=k=w=�=>>'>,>Q>�>�>�>??:?�?    @   000I0�0�0�011C1�1�1�1�12,2�4�49 9*9S;`;�;�;�?�?�?     �   40G0g0z0�0�0�0�011/1K1^1x1�1�1�1�1�1�12C2R2�2�233D3k3w3�344'4,4Q4�4�4�455:5
616G6e6�6�6�6727R7�7�7�78-8@8D8H8L8]8b8l8�8�8�8�8�8S9`9�9:�:�:�:�:�:�:�:#;1;�;�;�;<=+=A?e?�?�?�?�?�? 0 |   000!0c0r0�0�2[5s566s6�6�67C8P8�8�8;9S9�9�9�9�9Y:k:�:�:�;�;I<[<�<�<=+=c=s=�=�=>'>0>8>�>�>�>??R?�?�?�?�?�?�?�? @ �   000&0-0;0F0_00�0�0�0111f1o1v1}1�1�1�1�122D2�2�2�2�2�2�234�5�5�5�56>6G6P6X6�6�6�67$7S8`8�8�8< <�<�<�<*=�=�=�>�>{?�?�?�? P @   $0y0�0O12I2w2�2�2�4�4%6+686A6J6S6,9t9e:3;�>�>?0?�?�?�? ` H   �01181=11�1�1�1"2'2I2V2y2~2�243s3�3�3�3�3�3�3�344#4.4O4)>;> p 4   30E0D13.3�3�34%4;4I7Q7H8p:x:�;�;�<>>^?�?�? � H   {0�0�0�0�0�0�0j34u4w6�6�67777"7+7;7C7�7;8]8l819a<�<B=d=�=   �    t0�0�0C3T334F4�<'>W? �    �4�4�9:r;�?�?   � l   33]3f3o3w3�3�3�4O6X6a6i6r66B7K7T7\7e7n7�788�8 9'979�:s;�;�;�;< <c<p<�<�<=3=C=l=�=>�>?"?�?�? � @   0,0�083L3�4�4�8�8S=c=�=�=�=�=�=�=>>*>u>�>�>????? � d   #404�4�4535j5�5�5�5�5�5�56)6[6n6}6�6�6�6�6�67*7=7D7W7r7�7�7#828�8�8�;�<�=�=�=D>I>S>�?�?   � P   �0�0�0�0�2�3�3D;I;S;�;�;�;�;�;�;<<<s<�<�<�<�=�=�=�=�=�=>J>q>�>�>:?a? � l   0(0M0r0�0�0�0
111"2L2}2�2�2�2�2�2�2373i3�3�3&4J4q4�4�4M6[6m6�6�6a7s7�7�7�7�89@9�99:�:�:�:�:�:�:     @   T3�3�3�4�4�9�9:3:�:�:[<s<�<�<d=o=�=�=�= >$>0>e>�>�>�?�?  �   0)0Z0�3�3�3�4�4Y5k5�6�6�6777u7�7�7�788s8�89{9�9:$:C:y:�:�:;2;L;�;�;	<#<�<�<�<�<$===`=t=�=�=�=>&>Z>s>�>�>	?"?�?�?�?     �   0@0]0{0�0�0�011F1�1&2D2n2�2�2�2�23^3s3�3�3�3�3�3484W4s4�4�4�4�455 5$5(5,5054585I5^5�5�56!6Y6x6�6�6�7�7838Y8t8�8�8�8999X9�9�9�:/;S;�;,<\<�<�<=�=�=�=�=>">�>�>F?_?v?�?�?�?�?�?   0 �   090U0l0�0�0�0�01)1L1s1�1�1�12(2Y2n2�253E4`4�4�4�4�45$5N5c5�56?6V6}6�6�6�6�67@7^7�7�7�7�7�7888�8�8�9�9�9
:;:Z:e:�:�:�:�:;3;R;�;�;
<U<�<�<9=K=�>? @ @   92M2�3�38�8�89999%9*949X9]9g9 ::::�:�:�:4<(=?   P �   )1=1�1`2
555]5b5l5)6;6�6�67#7H7[7�7�78$8=8c8s8�8�8�8�8999X9::K:^:�:�:�:�:#;3;h;{;�;<#<4<X<]<�<�<�<�<�<�<�<M=y=�=�=�= ` X   X0�1/444>4�4�4�4c5v5�6�6A7}7�7�7�7�7�7�708�8�8s9�9�9�9�9(:�:�:�:;-;Z;v;�;<C<   p d   l0�0�0�01$1C1b1�1�1�1�1�1292[2�2�2�2%8+8�8�9:+:Q:u:�:�:/;;;�;�;<4<T<{<�<�<�<=o=t=�?�?�? � P   !0`0�1�1�133[3�3�3�34Q4�4�4�4595Q5d5�5�5�5�5�5�5�5�5�;�;5<�=�=�=U?�?   � D   �1�1T3�3�3L4Q4[4c5v5$6)63637F7�7�78*9/999;�;�;=(=C=U=!?8? � 4   S0.1H1y1�1�1%2�2�2<3t4�4�4c598d8{8�8�8�;�;   � �   0"0N0T0b0�0�0�0�0�031C1y11�1#202�2�233@3�3�3C4V4�5�566�6�67"7Y9n9�9�9�9�9�9::#:5:G:W;�;�;�<==f=>v>�>?�?�?�?�?�? � �   b0�0�0�0�1!2c2�2�2�2�2�2�2~3�3�3�3�344)4:4P4n4�4�4�45555%5<5C5a5�5�5�5$6,666@6J6T6^6h6w6|6�6�6�6�6�6�6�6�6�6+89n9(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:�<�<=="=�=�=S>e>�>?   �    	22�2�3�5�6�78 � X   �011"141C1S1{1�1�1�1�1�12S2a2z2�2�2�2�2�2}3�3�3�3�3�3�3"4c4v4�48)8C;W;�=�=   � \   5%5G5�6�6L7Q7[7b8g8q8�8�8�9�9�9�:�:�:�:�:�:S;f;<<"<\=a=k=�=�=�=S>f>??"?�?�?�?     X   O0T0^0�0�0�1�1�1�1�1�1Y2^2h2*3/393�3�3�344�4`5�5�5	7�7�7�8�8�9�9�9�9�9:�?�?�?  p   0 0�0�01#1S1`1�1�1!2R2b2r2�2�2�23#464�5�5�67�8�8�8-9�9G:L:V:�:�:�;�;�<�<�<�<Z=�=�=�=�=�>�>?N?�?�?�?   D   C0R0�015122c2q2#515�5�5S6d67C7r7�7�<�<3=@=�=�=s>�>�?�?   0 h   �0�0�1�1�2�2c3p3�3�34474?4H4P4�6y7�7�8�9�9�9:F:s:�:�:+;�;�;�;A<s<�<=@=y=�=�=->�>�>�>E?w?�?   @ h   0C0|0�01T1�1�12e2�2�263h3�3
4�4�4�5�5�566!67�7�7�7R8W8a8�:�:�;�;`<�<P=w=@>g>�>>?P?�?�?�?�? P x    020�0�0�0�1�1�2�233E3�3�3?4�4�4S5�56�67G7L7R7_7�7�788j8�8�8�8�819C99:K:s:�:�:	;+;�;�<�<= =V=�=/>g>O?w?�?   ` P   	00�0�01+1i1{1�;�;<+<Y<k<�<�<�=�=>2>R>e>�>�>�>�>�>�>?!?>?Q?�?�?�?�? p t   �0�0�0S1X1�1�122 2b2�2�2$363E3�3�3�4�4�4�4575�566]6t6�6�6�6c7h7�7�78%8\8�8�8J9`9�9�9�9C:H:�:�:�:$<;<�< � @   0b0�12D3T3d3t34U4�4�4'5W5�6�6�6g:�:�:�:<< <c=u=�=   �     030E0W073c3u3�3s6�6@?   � p   ^0�1�1w2\3r3�344!455�7�78%8;8�8�8�9�9�9�;�;<7<e<�<�<�<�<�<==E=a=k=�=�=S>c>|>�>?=?T?{?�?�?�?�?�? � 8   0010y2�3�3�45c5r5�5C7U7g7�7B8�9�:H;b<b=�=?�? � �   �0R1[2�2P3�3�4�4�4�45)575\5j5�5�5�5�566�6�6#7�7�7�8�8�8�9�9:Z:�:�:�:�:�:;5;;�;�;
<$</<{<�<�<{=�=�=�=�=�=(>L>�>Y?�?�?�?�?�? � �   0*0~011a1f1q1�1�1�12V2393>3I3g3r3�3�304�455!5?5J5�5�56�6�6�6�67!7i7�7�7�8�8�8�8�8�8x9�9�9v:�:�:�:;;V;z;�;�<�<�<�<�<�<?=\={=*>Z>_>j>�>�>�> ?M?X?�?�?�?   � d   _0�0�0�0�0�0151]1h1�1�122,272�2�2�2�2�34?4�4}5U6#717Z7�7�7�7�:;;�;6<<<x<~<�<�<B?�?�?�?�? � �   �1�1�1�1�1�132@2�2�2�2[3s3�3�3�3�3444 4,434D4R4_4f4t44�4�45+5o5�5�5�5�5�5 6+6L6W6x6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�8Y9n9�9,:C::�:�:@<�<==== =$=(=,=0=A=R=�=J>q>�>�>�>?     �   u1�1�1�1�1C2L2U2]2�2�2�2�2^3j3u3�3�3�3�3(4,4044484<4@4D4�4�4�46666z6�6�6727G7_7d7t7�7�7�7�7�7�7�7�78808@8G8U8|8�8�8�8�8�8�8�8�9�97:?:G:P:�:;;(;7;^;�;�;<U<�<{=�>�>�>�>�>    d   .0f0�0�0Z1o1�1�2
3^3�3w4�4�455J5�516;6�89.9d9�9�9�9$:(:,:0:4:8:�:�;�;�;�;�;�;�;�;�?�?�?�?   d   00060A0Z0e0~0�0�0�0�0�0�0�0�011!101;1O1Z1v1�1k2�2�2�2�2+6C6s6�6�6S8f8�8r9�9�9t:�:u;#<6< 0 h   c0p0�0�0S1`1�1�1A2I2Q2Z2�6�6�6�6�6;9S9�9�9�9�9Y:e:p:|:�:�:�:@;G;�;�;�;�;�;�;�=�=�=>#?0?G?�?�?   @ d   90N0�0�8�89(9�9�9�92:7:>:�:�:�:n;�;�;�;�;�;�;�;<<<1<D<^<�<�<�<�<=\=�=�=�=>O>�>?d?z?   P �   0F0�0�01\1�1�1'2g2�2�2343}3�3�3g5�5K6�6B7W7�7�7�7�7�8�8�89B9[9�9�9:6:O:m:�:�:�:;l;�;�;�;
<<H<b<w<�<�<�<�<�< =	===#=,=4===F=N=W=`=k=w=�=�=�=�=�=�=�=�=�=(>S>_>k>v>�>�>�>�>�>�>�>�>
?�?   ` (   O2p2�2�4�;
<<+<2<@<y<=$=.=�?   p @   �0�0�0�1�1V2�2�3�3�3#404�4�4535e5#9(9291:6:@:Y=m=Y?m?   � �   �2�2*3_3�3y4�4�4�4�4�4�4�4�4�4�4�4555!5*535<5E5R5[5d5m5�5�5�5�5�5�5�5�5�5�5�5�5T6y67&7�781888?8Q8X8^8s8�8�8�8�8�8�8�89949?9X9c99�9�9�9::$:=:D:J:\:c:i:t:�:�:�:�:�:�:;;6;A;_;j;�;�;�;�;<< <<<N<`<r<�<�<�<�<�>�>?`?�?   � �   �2�2�2�2�2�2�2�2�2333#3-373A3K3U3_3i3s3}3�3�3�3�3�3�3�3�34.4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�455�5�5�56�6�67c7q7 � ,   �0�0J1J2�6�6�;�;�;�;
<�<a=f=p=C>R>a> � ,   #353G3x3~3�3�3�3�388�8�8�8�8�>�>? � |   �0�1`4d4h4l4p4t4x4|4�4�4�4�4�4�4H5L5P5T5X5\5`5d5h5l5p5�9�9�9�9;;;;.;7;@;I;R;c<q<�<�<=c=t=�=>>c>r>�>�?�?�?�?   � X   �0�0H1{1�1�1�1�1�2�2�2�2�2�2�2�2�23�3�3�3�3�3�3�3�3�3�3�3i;{;Y<k<�>�>�>�>?�?   � l   0�0�0�0�0�2�3	4k6�6�6�8�8�8�8�8�8�8�8�8�8�8999!9*939<9�9�9�9�9�:;";�;�;j<�<�<�=�=�=#?5?F?�?�?   � p   1 1$1(1,1D1�155�7�7�7�78 8*8l8p8t8x8|8�8�8�8�8�8�8�8�8�8�8�9m;{;�;=�=�=�=>>D>K>�>	??;?A?G?P?�?    	 �   i0{0191K1�1�1�1�1252;2A22�2�2�2�2�2O3m3�3�3�3�34-4H4{4�4�4�4�45A5R56[6j6�6�6�6�67�7�7�7�78"8y8�8�8�89"9�9�9::D:�:�:;w;�;<h<4=9=C=x=}=�=�=   	 �   �0�01101B1T1f1X2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,30343�5�8�8 91:C:S::�:�:�:�:�:;;*;u;.<3<=<�=�=�=!>&>0>? ?*?�?�?�?  	 (   �2�2�2�2�3�3R4j4495K5�5�6�6�6   0	 d   �0�0�0#131�1�1�2�2�2W3\3f3{3�3�3�3�34441464T4�5�5�8�8�8�8+9�9�9�9(:;:X:k:�:�:�:;;*;/;9; @	 $   =0B0L0�0�0�0�01�8D9�:�:�:   P	 \   �3�3�3k4p4~4�4�4�4=5B5s5x5�5666�8�8�8�9�9�9�;�;)<.<�<�<�<�<�<J=O=�=�=�=�>�>�>�?�? `	 d   000I2[2�2�2�2�2+303:3�3�3�3�3�3�4595>5H5�5�5�5,616�6�6�6�9�9:M:c:r:�:�:�:;0;�;S=e=S?e? p	 H   92_2�8�8�899�9�9�9c<h<r<�<�<�<�<�<�<h=m=w=�=�=�= >>>->2><>   �	 �   -066%6b6g6q6�6�6�6�677-727<7]7b7l7�7�7�7�7�7�7l8q8�8�8�8�8�8�8(9-9H9M9W9�9Z:|:�:�:�:�:�:�:�:�:�:T;�;�;1<6<@<_<�<�<�<�<;=@=J=C>H>R>�?�?�? �	 ,   C0V0�2�2�2�34,4�7�7�9�9�9;&;�>^?�? �	 @   x0_1�1�13$3G3�3 44!4y4�4�4�4�4�4788�9�9i;{;�;�;�?   �	 H   �0�0\1�3�5l7p7t7x7|7�7�7�7�7�7F9�;<	<B<G<Q<�<	??Y?^?�?�?�?�?�? �	     K0P0Z077C:V:�=�=�>�>�? �	     0�12�4�436I6~;�>�>�>�> �	 �   -121<1�1�1�1�1�1 233M3`3S4i4{4�7�7�7c8h8r8�8�8�8�9�9�9Q;n;s;};�;�;�;<<<<0<5<;<E<X<^<d<m<�=�=�=>>>>&>N>S>]>�>�>�>?	??0?5???]?b?l? �	 |   1$1z4�4�4�4�4�4�4�4�4%5*545N5S5]5w5|5�5�5�5�5�5�5�566 6�6�6�6�677"7'717`7e7o7�8�8�8�<�<�<�<�<�<�<n>s>}>�>�>�>    
 �   0D0�011B1a1�1�1�122?2D2N2d2i2s2d4�4�4�45#5-5i5n5x5�5�5�5�5&6+656z66�6�6�6�6�6�67*7/797^7c7m7�7<8A8K8{8�8�8!9&909�9:�:�:�:�:�:�:�:�:;�<�<�<,=1=;=s=y=�=�=�=�>?�?   
 �   0�0'1�192�2:3�3�3�3�355)5�5�5�5�5�5 6B6G6Q6t6y6�6�6�677*7/7978$8.899'9Q9V9`9�;�=�=�=H>L>P>T>X>\>`>y>~>�>+?0?:?�?�?�?  
 �   )0.080c0s0�0�0�0�0�0�0]2b2l2�2�2�2d3i3z33�3�3�3�3�3E4J4T4�4�4�4$5)5:5?5I5�5�5�5�5�56M6R6\6�6�6�6�6�6:7?7I7�7�7�7�788�8�8�8�8�8�8�8�8E9J9T9s9�9�9�9�9r:w:�:�:�:�:�:*;/;9;�;�;�;�;�;<�<�<�<�<�<�<�<�<U=Z=d=�=�=�=4>9>J>O>Y>�>�>�>???�?�?�?�?   0
 �   0M0R0\0�0�0�0�1�1�1�1�1�1�1�1W2\2f21363M3R3\3�3�3�3�4�45\5a5k5666w6|6�6772777A7k9p9z9P:U:_:�:�:�:@;�<�<d=p=�=�> ?$?(?,?0?4?8?<?@?D?H?L?P?T?X?\?`?d?h?l?p?t?x?|?�?�?   @
 �  0000F0�0�0�0�0�01$1.191D1O1Z1e1s1~1�1�1�1�1�1�1�1�122:2K2a2w2�2�2�2�2�2�2�2�2�2�23333'30393B3K3T3e3�3�3�3�3�3�3�3�3�34434I4_4u4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5054585<5@5D5H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5064686<6@6D6H6L6P6T6X6\6`6~6�6�6�6�6�6�6�6�6�6�6�6�6�67(7,70747�7�7�7�7�7�7 8888888818P8T8X8\8�8�8�8�8�8�8�8�889<9@9D9H9L9P9T9X9C;Q;j;<&<I<�<�<S=f=�=�=+>�>?�? P
 |   �0�0�0W1e1�1�1�122$2_2�2�2�2�2�23?3�3�34�4�4W5�5�5U6�6�6�6�6+7@7�7�7858t8�8�89C9g9�9�9:?:�:�:;!;=;F;�;�;!<Z? `
 <   �0!1b1�1�1�1�1Q2r2�2�23�3�35�5�6�6�7�7�8�8i9~9&<D? p
    �0�6�6�>�>   �
 @   *1�1�2�2�5�5;7S7�7�7�7�7�78828E8�8�8�8�8�<�<="=�=�=|> �
 (   �566�6�6�8Q99;?;N;W;`;i;�=�=   �
 �   S0a0c2q2�2�2c4q4�4�45�5�5�5	6668!8�8!9�9�9':,:<:J:[:e:o:�:�:�:�:�:�:�:�:�:;1;8;R;a;h;m;};�;�;�;�;�;<<<<-<G<Q<g<q<�<�<�<�<�<�<�<�<=!=7=A=Q=Z=d=�=�=�=> �
 @   2M2y2�2�2�2�233�3�34;4V4{4�45�5�5�7�7�9�9	<<�>?   �
 0   �1�1A2a244�7�8�8�8�8�<=�=�=�=>?.?   �
     �2�35&58K8c8�8�8�:�=�= �
 (   �0�0C5Y5�5<6i68�8�8M9�9�:�:=   �
 X   �1�3:4�5�6�6�6�6�62777A7i7n7x7�9 :c:r:�: ;c;q;�;�;<5<j<�<�<�<*=<==?Y?�?�?�?�?     4   	010�12�7�7�8�8999$9.979m9�9�;�;"<o<�<�<  H   �2�5�5�5�5�67*7�8�8'9E9�:�:�;�;�;<{<�<�<�<�<3=A=j=|=�=�=�?�?     P   0&0
212s2�2�2�2�2�2�2'3t3�3�35K5x5�5�56'6W6q6�677"7;7T7�7�7�78;�;y= 0 0   �4�4�4�436A6j6�6�677i8~8�8	::�;�>�>�?   @ H   0y1�1<3V3x5�5�5$6�7�8�8�8�8�8#989%:�;�;�<�<== =*=4===�=�=6?Q? P D   �0�0S1b1�1�1#212J2�2�2+303
444>4C4M4�4�6:789.9V9q9;i?~? ` <   �1C3[3�455-5�7�7)8@8c8�8*9Y9�95:Y:�:�:<<�<�<=   p ,   0�0F28~8�8B:,;3;�;�;�<�<�<�<"=)?;? � (   s1�1�1�1�3�3i7{7	99�:�:�?�?�?   � |   0"0J0V0�0�0�0�0s1�1�1�1�1�4r5�5�5�5(6�67;7C7J7U7_7}7�7�7�7888(828<8x8�8�8�89959@9F9L9U9_9i9�9:�:;�;�;�>�>   � (   �0�1�3�3H58s8�8�:�:';�<%=1?F?   � 0   �0�0�0�0�0�1�4�4)6>6�7�7S;`;�;�;�<�=�=*? �     �0�23e4y4�6�6�6�6i9~9   � 4   81f3N4Y5n5�5�5t6�7
8v8�8�8�=�=>>>>p>�>�>�? � �   �0�0111H1Z1�1R2h2�2�2�2�254:4D4%6W6C7V7*8Q8c8r8�8�8�8�8�8�8�8�8�8�9:!:9:�:�:�:�:�:�:�:�:K;e;�;�;�;<]<�<�<�<�<�<�<=1>9>B>K>S>_>k>v>�>�>$?;?�?�?�? � |   S0b0�0�0C2Q2�2�2�34*4Q4#505�5�5�5K6c6�6�677*7�7�7L839l9r9�9�9C:Q:�:�:�:�:+;C;u;�;�;�=>3>C>c>q>�>�>�>�>�>�>??�?        0c0r0�1�6i7q:e;j<�<�<??     @1r2   l   �2�23/3Z3�34!4-484Y46!6�6�6�67%717<7H7S7_7919J9q9�9�9�9�9
:1:J:q:�:�:*;Q;c;s;%=-=O=W=}=�=�=�?   0 �   b1�1�1�1�12&2/282@2�3�3�3�3�3�45#5-5�5�5�56666'606S6�6�6�6727K7�8�899�9�9�9�9�9�9::5:[:s:�:�:�:�:;;!;);e;�;�;�;�;<.<O<X<a<i<�<�<�=�=+>C>�>�>�>�>#?0?�?�?   @ T   030�0�01k1�1�1�1F2a2w2�2�2�2�2�2A3G3�4K6�6�6�7�8]:�:�:�:�:i<�=�= >E>�>�>? P p   �0�0#2v2�2�2I3^3�3�344B5Y6�6�6#707�7�7+8C8�8�8�8+9t9�9:X:�:;;@;�;�;�;�;<B<i<~<�<=c=k=�=�=�=#>+>   ` x   1)1N1�1�1�2�2M3�3	4.4s4�4�4�4{5�5�5�5#626 77C7P7�7�738@8�8�8+9C9�9�9::O:b:&;2;;;D;M;V;s;�;=>>>>>)>>>�? p T   0�0�0;1R1�1�1v3�3	44�4�4)5>5s6�6)9>9X:p:�:�:�;�;2<�<�<�<�=�=F>]>�>�>�?�?   � `   i0{0141�1�1�1S2f293d3�4�4 5555.5	7�8�8#939Q9l9y9U:�:;+;;;<3<C<p<�<e=3>C>f>v>0?e?   � �   U0�0�0�0#121�1�12"2�2�233�3�3�3#424m4�4�4�4#525m5�5�5#626�67)7"8�8�8�8999K9�9�9�9�9	::S:d:}:�:�:;=;k;<&<H<j<�=�=�=>?!?,?Q?l?s?z?�? � X   b0�122�2�2�6�68>8h8o8�8�89}9�9(:�:�:;Y;�;�;�;&<Z<�<�<�<�<�<�<==�?�?�?�?   � @  �01R1[1s1�1�1�1�1�1�12252C2R2�2�2�2�2�2�2�2 3#313N3e3s3�3�3�3�3�3�34!404S4a4~4�4�4�4�4�455,5>5Q5`5�5�5�5�5�5�56636C6\6n6�6�6�6�6�6�677B7K7c7s7�7�7�7�7�7�78%838B8r8{8�8�8�8�8�8�89!9>9U9c9r9�9�9�9�9�9�9: :C:Q:n:�:�:�:S;b;�;�;�;�;�;�;�;�;�;�;#<4<M<�<�<==<=�=�=�=7>J>s>�>�>�>�>�>�>???#?P?`?�?�?�?   � x    00@0d0z0s2�233�3�3#414�4�4C5Q5�5�5c6q6�6�6K8+9�9R;[;s;�;�;�;<<#<1<J<`<�<�<;=S=�=�=�=�=�>�>�>??c?q?�?�?�? � h   31A1�1�1�2�2d3�3"4+4C4R4k4�4�4�4 66666666 6$6(6,60699c9q9�9�9�9�:�:;�<A=S=e=�=�=Y>�>�? � �   f0}0�0�0�0�0�0K1c1�1�1�1�12222.2:2E2Q2�2�3�3"4F4_4�4�4�4�56u6�68�8�8�89C9P9�9�9m:�:�:�:�:�:;3;J;g;�;�;�;�;�;�;�;�;�;'<C<R<y<�<�<�<�<i=|=�=�=�>�>?:?J?W?`?i?r?�? � �   �0�0�0�0-1>1�2�2�23
33)3A34 4�4�4)6@6W6�6�6�6�67)7U7h7|7�7�7�7i9|9�9�93:�:�:+;C;�;�;G<{<�<�<�<�<
===$=>=c=q=�=�=s?�?�?�?     h   �0�0�0�011*1c2p2�233�3�3#404<4Z4�4T5Z5y55�5I9[9�9�9�:;I;[;�<�<�<�<�<
=c=t=�=�=�=>>S>a>�>  <   C0P0�0�0�0�1�1M334g45�5�5�5�5�7�7�8�8::�:�:�?�?     p   0!0�0m1�1�1b4�4�4�4�4 555(5�5P6T6X6\6`6d6�7�7�7�7�7S:a:�:�:�:;{;�;�;<<A<�<�<�<=	=#=(=C?Q?j?o?�?   0 $   E0G3O3#535y9�9�;�;<!<y>�>   @ l   �1�1212A2F2P24!4�6�6�6�6�67!7s7�7�7�8.949:9E9Y:v:�:�:�:;!;:;3=@=�=�=�=[>s>�>�>?3?�?�?�?�?�?�?�? P h   C1T1�12C5R5�5�5�56&6@6�6�6�6�6�6 77Z7�7�7�7�788�8�8C:S:�:;�;�;=3=`=}=�=�=�=�=�=�=	>>�>   ` (   L0o1�6�6j7Q:3;B;�;<�<I=^=�=/>E> p (   �0_1�1L3P3T3X3\3)6>6j9�9�9:�<�< � P   h5l5p5t5x5|5�5�5�5�5�566�67Q7e7�7�89S9c9�9�:�:C;R;�;�;<#<<<�<�<�<!= � �   c0r0�0�0�0�02$2F2q22�2�2�3�3�34,4F4Y4s4�4�4�4�45{5�5�56*6Q6j6�6�6�6�67*7Q718U819S9a9�9�9C:Q:w::;a;s;�;�;�;�;�;X<�<�<�=�=�=�=>�>?"?;? � �   1Q1�1�1�1�1�1�1�2�2S3b3�34c4p4�4�4[5s5�5 6C6R6y6�6�6�67O7b79�9�9�9�9::k:�:�:�:�:#;2;K;K<j<�<�<�<�<�<===�=�=�=�=>3>B>}>�>�>?!?`?�?�?�?   � L   ;0S0�0�011�1�122H2c2r2�2�23e3�3�34J4q4�4�4549�9�9�< =C=P=�=? � H   00*0�3�3�3+4Z4a4s4�4�4�4<5�5�5�5�56j7o7�7�7�7e8j8t8r=w=�=�=   � P   A0F0O0T0]0b0k0p0y0~0�0�0�0�0�0�5�56#6[6�89C9R9y9�9�9:c:q:�:�:c<p<�<�< � L   
111C1Q1z1�1�1�155�5�5#626�6�677>7�7�7�78C8Q8j8�:; ;9;R;m;=m= � @   �3y4�438@8�8�8+9C9�9�9;;4;_;z;;�;�;�;�>�>�>�>??D?     @   �0�0�0�1�1�23�4�4�4Q5�5�5�6�67,7�8�8�<�<s=�=�>�>�?�?    8   M1Y1�2�2o4�56)7>7�:�:�;<==z=�=�=+>C>�>�>�?     4   0�4�4�5�5�5.6D6�8�8�9�9:�:�:�:;;;5;�=�= 0 T   A0F0P0s0�0�0�0191�1�1$6�697�8�8�8�8�89C9T99�9�9$:�:�:�:|=�=>>;>V>|>�>�> @ <   �1�133[3�395N56�6�6�8�9:; ;�;�;�;;<S<�<y=�=?�? P P   0.0�1;2�2�2I6]6�7�7�78P8�8�8�89c9�9�9&:g:c;�;�;�;�;<?<]<q<�=�=P>�>   ` T   .0F0�0�0�01i1~1�12}2�4�6777h7�7�7�7�7�7�8�8�9�9�:�:<<H<j<�<�<�<==+= p h   11'10191B1U1�1�1#26233j3�3�3�3�3G4T5}5�5�5�5�6�6D7Q7]7l7{7�7�7�7�89s9�9�9�93;8;B;s;�;�;�;a< � |   �0
111C1Q1j1�1
2292^2�2�2�2#303<3�6�6�7�7�78*8�8�8�89-9N9W9`9h9�9�9�9�9�9:::C:S:l:�:�:�:�:C;R;�;�;< <�<�<1=I= � X   1A1Z1�1�1�1*2Q2c2q2�2�2�2
3a3y3�3�3�3�4�4�4�4�:�:&;+;5;�;�=�=�=>">V>?#?S?b?�? � `   e1�1�1S4a4z4�4�4�4K5c5�5�5�5+6C6�6�627�7�7�7898W8u8�8�8F9[9t9�9�9�9�9�9!:�>�>	??]?�?�? � (   1!1<1L1�4�4�4�6�6�9;;; ;<<!? � (   0)0C2V2Y3n3�9�9c;v;�<�<J>�>]?   �    �1�1�1�1�2�2�2�6�6e7 � $   g4m4�4�4.646|6x7�:�:�:�:�;< �     �3�7�;�;�;�;r<�<=m?�?�?   D   1�1�1�1'3.3<3�5�567;7B7�8�89w;�;�;�;�<�<�>�>�>�>�>�?�?�?    X   p0�0�0�1�1 3%3/3F3K3U3�3�3�3�3�3�3V6]6g6�7�7�7S8X8b8�8�8�80979r9y9�9+;0;0=5=?=�?      �0�7�7�8 0    (;/;;;   @ �   b0�5�7�7�7�7�7�7�7�7�7�7�7�7888#8-868@8J8S8]8g8p8�8�8�8�8�8�8�8�8�8�8�8�8c9i9n9x9~9�9�9�9�9s:�:�:�:j;y;�;�;�<�<=s=�=�=>->s>�>   P `   W0�0�0M1a1�1�1�2�2�2#333�34(4	55�5�6�6�637D7�7�7�7�8�8k9q9�:�:.;<;�;�;< <s<�<,==�>   ` ,   +1s1�1�12�3�3L5�7 9&9�<�<�<�?�?�?   p �   0@0D0H0L0P0T0�0�0�2�2�2!3U3`3l3�3�374�4�4�4�4�4�4�4�4�4�4�4�4�4�4 555551589=9G9q9~9�9�9�9�9�9�9�9�9':�:�:�;<F<K<k<t<�=�=�=�=�=�=�=�=�=�=�=�=>M>y>�>�>�>�>�>�>�>�>�>�? � l   0;0N0\0�0�0�3�34�5�5�5�5�5�5�56c6q6i7~7�7�7�7�7�7�7�7z8�839;9�9;;;;a<s<�<�<�<�<�<�<�<�>�?�?   � X   �2�2+3C3~3�56&6�6�6l8�89�;�;�;�;�;�;�;�;�;�;�;�;�;�;p<�>�>�>�> ????"?.?3?   � 0   0#0f0k0�0M2R24�7�7�7�7�9�9;%;�<�<	=�? � @   <0@0D0H031E1T1�2355555 5$5(5,50545853;I;�>�>�>?   � 0   �1�1�1�2�2�2�2�2�2+606:6q6�6�6|;�;�;#>6> � 4   !454Q4�5�78=8s8�8�9:E:�:�:�:k;�;�;�;<�>�> � X   �12"2-2s2�2�2�2�23c5p5�5�5#626�6�7�7�9:e<C=Q=u=�=�>�>?/?O?e?�?�?�?�?�?�?�?   �    c0p0�0�0k1�1�8     T   �1�1=3]3Q5�5::5;:;D;�;�;�;�;<<�<�<�<o=t=~=???8?=?W?\?f?�?�?�?�?�?�?    X   a0f0p02171A1�1�1�12$2.2S2X2�4�4�4!6M6~6�6�8�8�8s9x9�9�9�9::�<�<�<?	??E?J?T?   H   �0�0�0�0�0�0�0�011�1�1,252>2F2s4�4�45"5�5�5�8�8�8�8�9e?�?�?   0     ?1g2v2�2�2O9u9�9/=U=d=   @ 0   1!1�2�3�3�5�6	7]7�7�7<c=�=�=�=6>k?�?�? P `   0�2�2�2 3!5�6K7 9d9�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;; ;$;(;,;0;4;8;<;@;D;H;L;P;T;   `    <9�:d;s;�;<�<�< p l   �0�0�0�3�3�3�3�8�8�89909:9T9^9p9z9�9�9�9�9�9�9�9�9:
::":6:@:L:Y:s:z:�:�:�:�:�:�:�:;;;A;�?�?�? � �   2$2/2=2)535P5[5h5r5�5�5>7O7W7^7c7k7�7�7�7839K9P9�;�;�;<%<r<�<�< =======#=)=-=2=8=<=B=F=L=P=V=Z=o=�=�=>>/>?)?�?�?�?�?�?   �    0Y0�0�0J11�1�1�1�1�1�1�12!2(2,2024282<2@2D2�2�2�2�2�233,33383<3@3a3�3�3�3�3�3�3�3�3�3�3*4044484<4�4�45(5/575<5@5D5m5�5�5�5�5�5�5�5�5�5�56$6(6,606�6�6�6�6�6�6�6�67M7T7X7\7`7d7h7l7p7�7�7�7�7�7b8~8B9�9::G:W:d:O;�;�;v<�<�<�<�<�<�< ===8===G={=�=�=�=�=�=>=>Y>q>�>�>X?c?�?�?   � �   "0'0<0�0�0�0�01J1X1�1�1�12222r2�23+3N3Y3k3�3�3E4W4�4�4�4�45y5�5�5�5�5�5�56B6�6�6�6�677727z7�7818:8B8b8�8	99%9G9]9o9�9�9-:G:T:�:�:�:�:�:�:�:�>�>	??   � l   ~1�2I3^3�3�3�3J4}4�4 5&5w5}5�5�5�5�5
6Q6e6�6�6�677'7�7�7�8�8�899R9�9�9�9�9: :2:@:�:�;R<�<i=�=? � <   �0�122>2�2�3�4�6�8�9<0<<<c<p<u<�<�<[=f=s=�=�=+>B> � �   ]0d01�89A9�9�9":j:�:;;%;.;A;K;R;Y;c;j;r;�;<7<D<t<�<�<�<c=�=�=�=�=�=�=>�>�>�>�>�>�>�>�>??!?;?E?[?e?�?�?�?�?�?�?�?�?�? � �   0�0�0C1N1X1]1m1�1�1�1�1�1�1�1�1�1�1�1�1�1�1y2�2�2�3�3�3�3�34G4M4T4�4�4�4�4�4�4 565?5K5�5�5
6q7�7�7�7�7�7�7�7)818;8T8^8q8�8�8�89�9�9�9I:h:�:�:�:;);1;9;P;i;�;�;�;�;�;�;�;<< <@<E<=(=�=?   � �    0I0�1d3y6�6�6�6�8�9�9::":.:C:I:]:d:�:�:�:�:�:�:�:�:�:�:;; ;&;/;;;I;O;[;a;n;x;~;�;�;�;�;�;�;�;.<4<^<d<�<�<�<(=K=U=�=�=�=�=�=>>>>0>>>E>K>a>f>n>t>{>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>???)?.?9?>?K?Y?_?o?�?�?�?�?   p   0!0K0V0�0�0�0�0�0�0�0�0�0�0�0�01111)12171=1G1P1[1g1l1|1�1�1�1�1�1�4�4 5r:+;�<==H=N=W=^=�= >�>?�?  �   �0�0�011&151P1q1�1�1�2�2&444W4�4�45#575l5�5�5�5�5�5�56696[6�6�6�6�6�6737;7l7u7�7�7�7�7�7�78!8-8C8L8U8�89>9R9�9�9�9�9�9:�:.;?;o;w;�;�;<(<1<<<<�<=K=R=�=�=�=I>�>�>'?�?�?�?�?     T   0W0�1�1�1�1�2�23a3�3�3�3�3!4�45n5y5�567 7�7>8V8�8�8�899�;h<�=�=�=`?   0 �   �0�0�0�0�011	1'2`2t2�2�2�233X3b3�3�3�34&4x4~4�4�4�4�4�465>5�5�5�5�5�5�5�5�5�56	6@6�6�6�6�6�67 7%7�7�7�7�7�7�7�7888)828>8G8N8X8^8d8�8�899"9�9:O:3;;;T;n;�;�; <<<!<)<5<Y<a<o<v<�<�<�<�<�<�<�<== =3=W=�=
>> >'>4>;>A>I>O>[>`> @ �   �0�0�0�0�0�0�0�011)141:1@1E1N1k1q1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�12"2(292�246@6s6�6�67�8�8�899b9j9v9�9�9::8:�:�:�:;!;1;=;F;�;�;�;><K<W<�<�<�<�<=6>>>F>�>�>�>T?a?�?�?�?�? P (  �0�0�0�0�0�0Y1e1m1y1�1�1222F2h2�3�3�3�3Y4e4u4�4�4�4�4�4#5/5�5	66%616N6T6i6�6�6�6Z7p7�7�7�7�7C8x8�8�8�8�8�8�899'949Z9u9|9�9�9�9�9�9�9�9�9�9::: :$:(:,:0:4:8:<:@:D:W:�:J;R;f;p;�;�;�;�;�;�;<< <,<8<D<P<�<�<�<�<�<�<�< ==$=0=<=t=�=�=�=�=�=�=�=�=I>Q>Y>a>>�>�>�>	??!?x?�?�?�?�?�?�?   ` @   �0�0L1�1�1�122+2(3n3v3�3�3�3 4%;i<�<�<v=�=�=�=!?<?�?   p |   10;0]0s182^2�2�223v3�3�34>4k4z4�4�4�4�4�4�45�5Y6|6�6�7O9e9s9�9�9�9�9:j:~:�:�:,;7;d;o;w;�;�;+<8<b<�<�<�<v>�>?Z?   � �   �0�1�1S2b2�2�2�3�3g4�4�45�5�5�5�5�5�5�5�566.6J6\6j6{6�6�6�6�6�67:7�8�8�899N9Z9{9�9�9:	;;H;O;x;�;�;�;�;<"<=<F<N<;=�=�=�=�=>>>,>8>C>n>�>`? � p   %0�0181C1w1�1�1�1�1�1�1�1Y2e2q3�3b5v5�5�56M6�6�6�6�67178828J8�8�8o9�9:�:Q;t;�;�<r=">I>\>�>�>)?]?�? � P   010Y0�0�0�1�1�1�1�1)2+3�3�4�5�5�5G879c:�:�:"<�=�=�=�=�=�=�=�=>)>�?�?   � |   M0�01�476R6h6~6�6�6�7]8�8�829�9�9�9$:1:?:o:�:;%;�;�;�;�;�;<<�<�<�<�<�<�< =J=R=o==�=�=�>�>�>�>�>?p?u?z??�?�?�? � d   00Y0^0e0j0q0v0�0�0�0z1�1�1�1�1�1�1�1�1�12F2�6�6�6�6777$7T7�7b8�8E9Q9�9�9�9�:�:�:b;�=�? � `   O0�041M1d1j1z11�1�1�1�1�1�1�1�1222-2�2�2�22494?4/5�5�5�67�8K9c9�9�9::8:�<�=�>�>�> � t   z0222"2&2*2.222�3�3�34)4;4M4_4q4�475T5~5�5�5�6�607J7P7c7p7x7�7�7�7�88;�;.<;<W<o<|<�<�<�<l>�>�>�>??7?   � T   �0�0�1U3c3k3x3�3�3�3�3�3�3�3�34�45A5e5�5�5n6�9�:�:a;C<�<�<�=�=�=:>Q>�>�?�?   H   �0�12$2�2�2�2|3�3�3N4757J:N:R:V:Z:^:b:f:j:n:r:v:�:W;o;~;�;	<.<  4   �5�9�9.:5:�:�:;@;�;_<x<~<�<�<�<�<�=�=,>�?     P   v0�0+151<1_1�1�23C3p3�3�4�425�5�5�56�;�;�;�;<:<j<�<�<�<\=>�>�>C?t?�? 0 �   1151?1�1�1232c2�2�2�233+3Z3�3�3�34J4z4�4�4�5�5�5�56!6)6@6Q6Y6p6�6�6�6-7h7�7�78=8m8�8�89C9j9�97:]:�:�:�:*;Z;�;�;#<J<z<�<�<=M=z=�=�=>:>�>�>�>
?:?s?�?�?�?   @ �   30Z0�0�0�091�1�12d2�2�2 3J3}3�3�3�34[4�4�4�45M5}5�5�56=6s6�6�6 7X7�7�7
8=8m8�8�8
9N9�9�98:�:�:(;c;�;�;/<G<�<�<O=g=�=�=8>j>�>�>?M?}?�?�? P �   0:0�0U1z1�1�162]2�2�2�2(3]3�3�34n4�4�45S5�5�56*6n6�67C7s7�7�788-9Z9�9�9�9:M:�:�:;t;�;�;*<Z<�<�<�<0=k=�=�=
>:>�>�>�>?P??�?�?   ` �   
0M0�0�0�01J1z1�1�122c2�2�2�23M3}3�3�34=4m45C5s5�5�5�5�6#7R7�7�7T8�8�8�8
9:9j9�9�9:=:m:;*;Z;�;�;�;<M<z<�<�<
=C=s=�=�=>3>c>�>�>�>#?Z?�?�? p �   @0j0�0�0�0*1p1�1�12P2�2�2�2'3`3�4 6=6�67C7w7�8�8�89M9�9�9:C:u:�:�:�:-;];�;�;<[<�<�<�< =]=�=�=�=#>S>z>�>�>
?:?w?�?�? � |   #0�0�01X1�1�12C2�203k3�3�3�4a5�5�5+6Y6�6�6�637c7�7�7�78[8�8�8�89S9�9�9�92:{:�:&;	<X<�<�<=-=]=�=�=�=D>s>�> ?*?~? � �   0*0]0�01b1�1�1
2�2�23B3j3�3�34u4�4�4
5E5�5�5�5A6u6�6�67^7�7�7
8K8z8�8�829Z9�9�9�9":J:�:�:#;M;};�;�;
<V<�<�<=*=j=�=�=�=5>e>�>�>�>K?z?�? � �   0w0�01I1�1�1�12M2�2�2k3�34I4�4�4�4"5�5�56P6z6�6�6D7�7�7 8-8]8�89�9:b:�:�:;:;j;�;�;�;-<]<�<�<�<8=j=�=�=>*>Z>�>�>�>%?J?�?�?�? � �   0M0�0�0�01C1p1�1�1�1-2]2�2�2�2A3j3�3�34J4�4�4�4*5Z5�5�5!6R6�6�6�67J7}7�7�78=8m8�8�8�8-9]9�9�9 :-:]:�:�:;:;j;�;�;�;*<Z<�<�<�<=J=z=�=�=
>E>�>�>�>?M?}?�?�? � �   0=0m0�0�0�0-1Z1�1�1�12U2z2�2�2
3=3m3�3�3
4C4m4�4�4�455p5�5�5�5*6]6�6�6�6�6.7Z7�7�7�7-8k8�8�8�8$9M9t9�9�9:h:�:�:(;Z;�;�;�;-<]<�<�<�<�<a=�=�=�=>J>�>�>�>-?]?�?�?   � �   #0J0z0�0�01q1�12=2j2�2�23*3]3�3�3�3O4�4�45M5}5�5�56=6m6�6�6�637]7�7�78J8�8�89M9�9�9�9:P:�:�:5;];�;�;<P<�<�<�<+=Z=�=�=�=>[>�>�>?T?z?�?�?   � �   0:0�0�01:1{1�1�1#2U2�2�2�293�3�3�3-4y4�4>5s5�56C6r6�6�6�6;7r7�7�7�7-8�8�889j9�9�9�9-:e:�:�:�:;M;z;�;�;<=<m<�<�<=:=p=�=�=�=*>Z>�>�>?:?~?�? � �   0*0h0�0�01g1�1�12M2}2�2�23=3j3�3�3"4R4�4�4W5�5�5�56M6�6�6�67=7s7�7�7
8=8m8�8;9u9�9�9:@:c:~:�:�:�: ;;-;M;o;�;�;�;�;�;�;�;�;�;<<!<1<6<;<@<E<J<T<a<f<k<p<u<z<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<======$=1=:=?=D=N=a=f=k=p=u=z=�=�=�=�=�=�=�=�=�=�=�=�=>>>>>>$>1>6>;>@>E>J>T>a>f>k>p>u>z>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ??
??!?&?+?0?5?:?D?Q?V?[?`?e?j?t?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   �  0000 0%0*040A0F0K0P0U0Z0d0q0v0{0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0111111$11161;1@1E1J1T1b1m1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12222 2%2*242B2N2T2^2{2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23333 3%3*343�3�3�3�3�3�3�3c4o4y4�4�4�4�4#5/595C5M5Z5d5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�56666 6%6*646A6F6K6P6U6Z6d6q6z66�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6777777$7:7Z7`7m7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7888 8%8*848A8F8K8P8U8Z8d8q8v8{8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8999999$91969;9@9E9J9T9a9f9k9p9u9z9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 ::
::!:&:+:0:5:::D:Q:V:[:`:e:j:t:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;; ;%;*;4;A;F;K;P;U;Z;d;q;v;{;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;
<!<&<+<0<5<:<D<Q<Z<_<d<n<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<==== =%=*=4=A=F=K=P=U=Z=d=q=v={=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>>>$>1>6>;>@>E>J>T>a>f>k>p>u>z>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ??
??!?(?-?2?7?A?Q?Z?_?d?n?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?  d  0000$0.0A0F0K0P0U0Z0d0q0v0{0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0111111$11161;1@1E1J1T1a1f1k1p1u1z1�1�1�1�1�1�1�1�1�1�1�1�1�123282=2B2G2L2Q2V2[2`2e2q2�2�2�2�2�2�23!313A3Q3a3q3�3�3�3�3�3�3�3�344!414A4Q4a4q4�4�4�4�455!515A5Q5a5�5�5�5�5�5�5�5�566!616A6Q6a6q6�6�6�6�6�6�6�6�677!717A7Q7a7q7�7�7�7�7�7�7�7�788!818A8Q8a8q8�8�8�8�8�8�8   l  l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,2024282<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3P3T3X3\3`3l3p3�3�3�3�3�3�3�3�3�3p4t4x4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5054585�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�6�6�6�6�6�688 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8�8�8�8:: :$:�:�:�:�:�;�;�;�;�;0<4<8<<<@<D<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$=(=,=0=4=8=<=@=D=H=L=P=T=X=\=`=d=h=l=�=�=�=�=�>�>�>�>�>�>�>H?L?P?T?X?\?   0 �   �0�0�0�0�0�0�0�0�0�0�0�0�0�0$6(6,6064686<6@6D6H6L6P6T6X6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 88888888 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8d8h8l8p8t8x8|8�8�8�8�8L:P:T:X:\:`:d:h:l:p:L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;   @ d  �0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 11111111 1$1(1,1014181<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4�4�4�4�4�4�4 5555064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7,7074787<7@7D7H7L7P7T7X7\7`7d7 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99999999 9$9(9,9094989<9@9D9H9L9P9T9X9\9`9d9h9l9p9t9x9|9�9�9�9�9�:�:�:�:�:�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<   P �   P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�40:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�; <<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ` �   014181<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22�5�5�5�5�5�5 66666666 6$6(6L7P7T7X7\7P=T=X=\=`=d=h=l=p=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=`?d?h?l?p?   � �  �8�8�8�8�8�8�8 99999999 9$9(9,9094989<9@9D9H9L9P9T9X9\9�9�9�9�9�9�9�9�9�9�9�9�9 :::::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;; ;$;(;,;0;4;8;<;@;D;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<   � �  666666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7�;�;�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<d=h=l=p=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>>>>>> >$>(>,>0>4>8><>@>D>H>L>P>T>X>\>`>d>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�> � �   024282<2@2p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5054585<5@5D5H5L5   � P   �;�;�;�;�;�;�;�;�;�;�;�;�;�;<< <$<(<,<0<4<8<<<@<D<H<L<P<T<�>�>�>�>�>   �   ,0004080<0@0D0H0L0P0T0X0\0`0d0h0l0p0t0�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�9�9�9�9�9�9 :::::::: :$:(:,:0:4:>>> >$>(>,>0>4>8><>@>D>H>L>P>T>X>\>`>d>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�? � P   h1l1p1t1x1|3�3�3�3�3�3�3�3�3�3(7,7074787<7@7D7H7L7P7T7X7\7`7d7h7l7p7t7     �   P7T7X7\7H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$<(<   0 X  �0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 11111111 1$1(1,1014181<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3P4T4X4\4`4d4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5054585<5@5D5H5L5P5T5X5\5`5d5h5l5p5t5�7�7�7�7�7�7�8�8�8�8�8�8�8�8�8�8 99999999 9$9(9,9094989<9@9D9H9L9P9T9X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? @ �  00 0$0(0,0004080<0@0D0H0L0P0T0X0@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�122 2$2(2,2024282<2@2D2H2L2P2T2X2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;; ;$;(;,;0;4;8;<;@;D;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$=(=,=0=4=8=<=@=D=H=L=P=T=X=\=`=d=h=l=p=t=x=|=�=�=�=�=�=�=�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>   P �  �1�1�1�1�1�1�1�1�1�1�1�1�1 2222224444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,60686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7(7,7074787<7@7D7H7L7P7T7X7\7`7d7h7l7p7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88888888 8$8(8,8084888<8@8D8H8 9$9(9,9094989<9@9D9H9L9P9T9X9\9`9d9h9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�;�;�;�;�;�;�;�;�;�;0=4=8=<=@=D=H=L=P=T=X=\=`=d=h=l=p=t=x=|=�=�=�=�=�=�=�=�>�>�>�>�>�>�>�>�>�>�>�>�>�>\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?   ` �   00000000 0$0(0,0004080<0@0D0H0L0P0T0X0\0`0d0h0l0p0t0x0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�081<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2222X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,60646H6L6P6T6X6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7`7d7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99P9T9X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;; ;$;(;,;0;4;8;<;@;D;H;L;P;T;X;\;`;d;h;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ????x?|?�?�?�? p �  �2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�46666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�7�7 88888888 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8d8h8l8p8t8x8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�88:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�=�=�=�= >>>>>>>> >$>(>,>0>4>8><>@>D>H>L>P>T>�>�>�>�>�>�>�>�>�>�>�>�>�>�>   �     0$0(0,0004080<0@0D0H0L0P0T0X0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,2024282<2@2D2H2L2P2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�4�4�4�4�4 55   � �   �7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7<;@;D;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <(<,<0<4<8<<<@<D<H<L<P<T<X<\<`<d<h<   � D   4181<1@1D1H1L1P1T1X1\1`1d1h1�1�1�1�1�1�1222(242@2L2X2d2   � 8   �7�7�7�7�7�7�7�7�7�79999 989<9@9p:t:x:|:�:�: � �   �3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55 � �  77�7�7�7�7�7�7�7�7�78888 8$8,8D8T8X8h8l8p8x8�8�8�8�8�8�8�8�8�8�899 9$9,9D9T9X9h9l9t9�9�9�9�9�9�9�9�9�9�9�9::,:0:@:D:L:d:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:;;;; ;(;@;P;T;d;h;l;p;x;�;�;�;�;�;�;�;�;�;�;�;�;�; << <0<4<D<H<L<P<X<p<�<�<�<�<�<�<�<�<�<�<�< ==== =8=H=L=\=`=h=�=�=�=�=�=�=�=�=�=�=�=�=�=>$>(>8><>D>\>l>p>�>�>�>�>�>�>�>�>�>�>�> ?????$?<?L?P?`?d?h?l?t?�?�?�?�?�?�?�?�?�?�?�? � �  00000@0D0T0X0`0x0�0�0�0�0�0�0�0�0�0�0�0�011 10141<1T1d1h1x1|1�1�1�1�1�1�1�1�1�1�1�1�122 2$282<2L2P2X2p2�2�2�2�2�2�2�2�2�2�2�2�2�2333,30343<3T3d3h3x3|3�3�3�3�3�3�3�3�3�3�3444,4<4@4P4T4X4`4x4�4�4�4�4�4�4�4�4�4�4�4�4�4 555$54585<5P5T5d5h5x5|5�5�5�5�5�5�5�5�5�5�5�56666 686H6L6\6`6d6h6p6�6�6�6�6�6�6�6�6�6�6�6�6 7777(787<7L7P7X7p7�7�7�7�7�7�7�7�7�7�7�7 888$8(808H8X8\8l8p8x8�8�8�8�8�8�8�8�8�8�8 99 90949D9H9P9h9x9|9�9�9�9�9�9�9�9�9�9�9::: :(:@:P:T:d:h:p:�:�:�:�:�:�:�:�:�:�:�:�: ;; ;0;4;D;H;L;P;X;p;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;< <$<4<8<@<X<h<l<|<�<�<�<�<�<�<�<�<�<�<�< ===== =(=@=P=T=d=h=l=p=t=|=�=�=�=�=�=�=�=�=�=�=�=�= >> >0>4>D>H>P>h>x>|>�>�>�>�>�>�>�>�>�>�>??? ?(?@?P?T?d?h?p?�?�?�?�?�?�?�?�?�?�?�?   � �   00(0,0<0@0H0`0p0t0�0�0�0�0�0�0�0�0�0�0�0�0�0 11(1,10141H1L1\1`1d1h1l1p1x1�1�1�1�1�1�1�1�1�1�1�1�1�1 2222(282<2L2P2T2X2`2x2�2�2�2�2�2�2�2�2�2�2�2�2�2 3333 3$34383<3D3\3l3p3�3�3�3�3�3�3�3�3�3�3�3�34444,4<4@4D4L4d4t4x4�4�4�4�4�4�4�4�4�4�4�4�4�4555(5,50545<5T5d5h5x5|5�5�5�5�5�5�5�5�5�5�5�5�56666 6$6,6D6T6X6h6l6|6�6�6�6�6�6�6�6�6�6�6�6 7777 787H7L7\7`7h7�7�7�7�7�7�7�7�7�7�7�7�78 8$84888@8X8h8l8|8�8�8�8�8�8�8�8�8�8�8�899909@9D9T9X9`9x9�9�9�9�9�9�9�9�9�9�9�9:::,:0:8:P:`:d:t:x:�:�:�:�:�:�:�:�:�:�:;;;(;8;<;L;P;X;p;�;�;�;�;�;�;�;�;�;�;�;�;<<<(<,<0<8<P<`<d<t<x<|<�<�<�<�<�<�<�<�<�<�<�<====4=D=H=X=\=`=h=�=�=�=�=�=�=�=�=�=�=�=�=�= >>(>,><>@>D>L>d>t>x>�>�>�>�>�>�>�>�>�>�>�>??? ?$?,?D?T?X?h?l?t?�?�?�?�?�?�?�?�?�?�?�?   �    000$04080H0L0P0T0\0t0�0�0�0�0�0�0�0�0�0�0�0111(1,141L1\1`1p1t1|1�1�1�1�1�1�1�1�1�1 222$24282H2L2P2X2p2�2�2�2�2�2�2�2�2�2�2�2�2�2333,30343<3T3d3h3x3|3�3�3�3�3�3�3�3�3�3�3�3444,40444<4T4X4p4�4�4�4�4�4�4�4�4�4�4�4�4 5555(585<5L5P5X5p5�5�5�5�5�5�5�5�5�5�5�5�5666(6,60686P6`6d6t6x6�6�6�6�6�6�6�6�6�6�6�6�6 777747D7H7X7\7`7d7h7p7�7�7�7�7�7�7�7�7�7�7�7�7 8888(888<8L8P8T8X8\8d8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�899,909@9D9T9X9\9`9h9�9�9�9�9�9�9�9�9�9�9�9�9�9 ::(:,:<:@:D:H:P:h:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;,;0;4;8;@;X;h;l;|;�;�;�;�;�;�;�;�;�;�;�;�;�;<<< <$<(<0<H<X<\<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�< ===== =$=,=D=T=X=h=l=p=t=x=�=�=�=�=�=�=�=�=�=�=�=�= >>>>> >(>@>P>T>d>h>p>�>�>�>�>�>�>�>�>�>�>�>�>??,?0?@?D?L?d?t?x?�?�?�?�?�?�?�?�?�?�? � (  0000$0<0L0P0`0d0l0�0�0�0�0�0�0�0�0�0�0�0�0 11(1,1<1@1D1L1d1t1x1�1�1�1�1�1�1�1�1�1�1�1�122 2$2(202H2X2\2l2p2t2|2�2�2�2�2�2�2�2�2�2�23333,3<3@3P3T3X3`3x3�3�3�3�3�3�3�3�3�3�3�3�3�34 4$44484<4D4\4l4p4�4�4�4�4�4�4�4�4�4�4�4�45555$5<5L5P5`5d5h5l5t5�5�5�5�5�5�5�5�5�5�5�5 666$64686H6L6T6l6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�677 70747D7H7L7P7T7\7t7�7�7�7�7�7�7�7�7�7�7�7�7�7�78888,8<8@8P8T8X8\8d8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99 90949D9H9L9P9X9p9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9:$:(:8:<:@:D:H:P:h:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:; ;$;4;8;<;@;D;L;d;t;x;�;�;�;�;�;�;�;�;�;�;�;�;<< <$<(<,<4<L<\<`<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�< ====(=,=0=4=8=@=X=h=l=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>(>,><>@>D>L>d>t>x>�>�>�>�>�>�>�>�>�>�>�>�> ???$?(?,?4?L?\?`?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?        00000 0(0@0P0T0d0h0p0�0�0�0�0�0�0�0�0�0�0�0 11(1,1<1@1D1H1P1h1x1|1�1�1�1�1�1�1�1�1�1�1�122 2$2,2D2T2X2h2l2p2x2�2�2�2�2�2�2�2�2�2�2 33333,3<3@3P3T3X3`3x3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44(4,4<4@4D4L4d4t4x4�4�4�4�4�4�4�4�4�4�4�4�455 5$54585<5D5\5  P  �3�3�3�3�3�3�34444$404P4X4`4h4p4x4�4�4�4�4�4�45555$5,545<5D5L5T5\5d5l5t5|5�5�5�5�5�5�5�5�5�5�5�5�5 66646<6D6H6P6d6l6�6�6�6�6�6�67777$7,747<7D7L7T7\7d7l7t7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78888$8,888X8`8h8t8�8�8�8�8�8�8�8�8�8�8 9999$9D9P9p9|9�9�9�9�9�9�9�9�9�9 :::: :(:0:8:@:H:P:X:`:h:p:x:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;; ;(;0;8;@;H;P;X;`;h;p;x;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<< <(<0<8<@<H<P<X<`<h<p<x<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ==== =(=0=8=@=H=P=X=`=h=p=x=�=�=�=�=�=�=�=�=�=�=>(><>D>P>p>|>�>�>�>�>�>�>�>�>�>?? ?,?L?X?x?�?�?�?�?�?�?     $  0000$0,040<0D0L0T0\0d0l0t0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01111$1,181X1d1�1�1�1�1�1�1�1�1�1�1�1�1 22,242<2H2l2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23333$3,343<3D3L3T3\3d3l3t3|3�3�3�3�3�3�3�3�3�3�3�3�3�34444@4`4l4�4�4�4�4�4�455<5D5L5X5x5|5�5�5�5�5�5�5�5�56(646T6`6�6�6�6�6�6�6�6�6�6 7777$7D7L7X7x7�7�7�7�7�7�78(848T8`8�8�8�8�8�8�8�8�8�89(9H9T9t9�9�9�9�9�9�9�9::4:@:`:l:�:�:�:�:�:�:�:�:;;;;$;,;8;X;d;�;�;�;�;�;�;<<4<@<`<h<p<|<�<�<�<�<�<�<==0=8=D=d=l=x=�=�=�=�=�=�=>(>H>T>t>|>�>�>�>�>�>�>�>??<?H?h?t?�?�?�?�?�?�?   0 �  0$0D0P0p0|0�0�0�0�0�0 1 1,1L1T1\1h1�1�1�1�1�1�1�1�1�12242<2D2L2X2x2�2�2�2�2�2�2�2�23 3@3L3l3x3�3�3�3�3�3�34(4H4T4t4�4�4�4�4�4�45$505P5\5|5�5�5�5�5�5 66,646@6`6l6�6�6�6�6�6�6�6�67707<7\7h7�7�7�7�7�7�7�78 8@8H8T8x8�8�8�8�8�8�8�8�8�8�8�8�8�8 99,949<9D9L9T9\9d9l9t9|9�9�9�9�9�9�9�9�9 :$:D:L:T:\:d:l:t:|:�:�:�:�:�:�:�:�:�:;;;;$;,;4;<;D;L;T;\;d;l;t;�;�;�;�;�;�; <<,<4<@<`<h<t<�<�<�<�<�<�<=$=D=P=p=|=�=�=�=�=�=�=�=�=�= >>>4><>D>L>T>\>d>l>t>|>�>�>�>�>�>�>�>�>? ?(?4?T?`?�?�?�?�?�?�?�? @ �  00 0@0L0l0t0|0�0�0�0�0�0�0�0�01 1(101<1\1h1�1�1�1�1�1�1�1�12$2,282X2d2�2�2�2�2�2�2�2343<3D3L3T3\3h3�3�3�3�3�3�34484@4H4P4\4�4�4�4�4�4�4�4�4�4�45555$5,545<5D5P5p5|5�5�5�5�5�5 6 6,6L6T6\6d6p6�6�6�6�6�6�6�6 7777$7D7P7p7|7�7�7�7�7�7�7880888D8d8p8�8�8�8�8�8�8�89$909P9\9|9�9�9�9�9�9�9�9�9: :,:L:T:`:�:�:�:�:�:�:�:�:�: ;;;4;@;d;�;�;�;�;�;�;�;�;�;�;�;< <@<L<l<x<�<�<�<�<�<�<�<=== =,=L=X=x=�=�=�=�=�=�=>(>4>T>`>�>�>�>�>�>�>??0?<?`?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   P �  0080D0d0p0�0�0�0�0�0�0�0 1111 1(141T1\1d1l1t1|1�1�1�1�1�1�1�1�1�1�1�1�12$2,242@2d2�2�2�2�2�2�2�2�2�2�2�23(3H3\3|3�3�3�3�3�3 4444$4D4P4p4|4�4�4�4�4�4�45555$5,545<5H5h5t5�5�5�5�5�5�56$6D6P6p6|6�6�6�6�6�6 7 7,7L7X7x7�7�7�7�7�7�78(848T8`8�8�8�8�8�8�8999 9@9L9p9�9�9�9�9�9�9�9�9�9�9:$:D:P:p:|:�:�:�:�:�: ; ;,;L;X;x;�;�;�;�;,<\<t<�<�<�<�<�<�<=$=,=4=<=D=L=T=\=d=l=t=|=�=�=�=�=�=�=�=�=�=�=�=�= >>>> >(>0>8>@>H>P>X>`>h>p>x>�>�>�>�>�>�>�>�>�>�>?,?4?<?D?L?T?\?d?p?�?�?�?�?�?�?�? ` �   0000 0(00080@0H0P0X0`0h0p0x0�0�0�0�0�0�0�011<1\1d1l1t1|1�1�1�1�1�1�1�1�1�12(202<2\2h2�2�2�2�2�2�23383D3d3p3�3�3�3�3�3�3�3�3�3�3 4 4,4L4X4x4�4�4�4�4�4�4�45585D5d5p5�5�5�5�5�5�56 6@6L6l6x6�6�6�6�6�6�67$7,787X7d7�7�7�7�7�7�7�7�7�7�7�7�78$8,888X8`8l8�8�8�8�8�8�8�8�89(949X9x9�9�9�9�9�9�9�9�9�9�9�9�9�9:::8:D:d:p:�:�:�:�:�:�:�:�:�:�:�:;;; ;@;H;P;X;`;h;p;x;�;�;�;�;�;�;�;�;�;�;<<4<@<`<l<�<�<�<�<�<�<�<=$=D=P=p=|=�=�=�=�=�=�=>(>0><>\>d>p>�>�>�>�>�>�>? ?@?L?l?t?�?�?�?�?�?�?�?�?�?�? p    00080@0L0p0�0�0�0�0�0�0�0�0�0�0�01111$1,141<1D1L1T1\1h1�1�1�1�1�1�1�1 22242@2`2l2�2�2�2�2�2�233 3(343T3`3�3�3�3�3�3�3�3�344(4L4l4t4|4�4�4�4�4�4�4�4�4�45,5L5T5\5d5l5t5|5�5�5�5�5�5�5�5�5�5�5666$6,646<6H6h6t6�6�6�6�6�6�6�6�6�6�6 77747@7`7h7t7�7�7�7�7�7�78$8H8h8p8x8�8�8�8�8�8�8�8�8�89$9,989X9`9h9p9|9�9�9�9�9�9�9:::8:@:L:l:x:�:�:�:�:�:�:�:;;; ;,;L;T;`;�;�;�;�;�;�;�;�;�;<(<H<P<\<|<�<�<�<�<�<�<�<�<=$=D=L=X=x=�=�=�=�=�=�=>(>0>8>@>H>P>X>`>h>t>�>�>�>�>�>�>?$?D?P?p?|?�?�?�?�?�?�? �    000080@0L0l0x0�0�0�0�0�0�0 11,181X1`1l1�1�1�1�1�1�1�1�12(242T2\2d2l2x2�2�2�2�2�2�2 3333<3D3L3T3`3�3�3�3�3�3�3�3�3�3 44444@4`4l4�4�4�4�4�4�4545<5D5L5T5\5d5l5t5�5�5�5�5�5�5�5�5�5 6 6(60686@6H6T6t6|6�6�6�6�6�6�6�6�67 7,7L7T7`7�7�7�7�7�7�7�7�7�7�7�7�7�7880888D8d8l8t8�8�8�8�8�8�8 99,949<9D9P9p9x9�9�9�9�9�9�9�9�9: :@:L:p:�:�:�:�:�:�:�:�:�:�:�:;(;0;8;@;H;P;X;`;h;t;�;�;�;�;�;�;�;�;�;�;�;�;�; < <(<0<<<\<d<l<x<�<�<�<�<�<�<=(=H=T=t=�=�=�=�=�=�=>$>0>P>\>|>�>�>�>�>�>�>??4?<?H?h?t?�?�?�?�?�?�? � �  0 0,0L0T0`0�0�0�0�0�0�0�01181D1d1p1�1�1�1�1�1�12 2@2L2l2x2�2�2�2�2�2�23(3H3T3t3�3�3�3�3�3�3 4444<4H4h4p4|4�4�4�4�4�4�45(505<5\5h5�5�5�5�5�5�5�566(6H6T6t6|6�6�6�6�6�6�6�6�6 7 7,7L7X7x7�7�7�7�7�7�78(848T8`8�8�8�8�8�8�89909<9\9h9�9�9�9�9�9�9:::(:H:T:t:�:�:�:�:�:�:�:�:�:;$;D;P;p;|;�;�;�;�;�; < <,<L<X<x<�<�<�<�<�<�<=(=4=T=`=�=�=�=�=�=�=>>>8>@>H>P>\>|>�>�>�>�>�> ??,?8?X?d?�?�?�?�?�?�? � �  0040@0`0l0�0�0�0�0�0�011<1H1h1t1�1�1�1�1�1�1 2 2,2L2X2x2�2�2�2�2�2�23(30383D3d3p3�3�3�3�3�3�34 4@4L4l4t4�4�4�4�4�4�4�45545@5`5l5�5�5�5�5�5�5�5 6 6(606<6\6h6�6�6�6�6�6�6�6�67(7H7T7t7�7�7�7�7�7�7 88848<8D8P8p8|8�8�8�8�8�8�8�8�8�89$9,949@9`9l9�9�9�9�9�9�9�9 : :,:L:X:x:�:�:�:�:�:�:�:�:;;(;L;l;t;|;�;�;�;�;�;�;�;�;�;<<0<<<\<h<�<�<�<�<�<�<�<�<=$=0=P=\=|=�=�=�=�=�=�=�=�=>$>D>P>p>|>�>�>�>�>�> ? ?(?0?8?@?H?P?\?�?�?�?�?�?�?�?�?�?�?   � �  0000<0\0h0�0�0�0�0�0�0�01 1@1L1l1x1�1�1�1�1�1�1�1222 2(202<2\2d2p2�2�2�2�2�2�23 3@3L3l3x3�3�3�3�3�3�34(4H4T4t4�4�4�4�4�4�45$5,545<5D5L5T5`5�5�5�5�5�5�5�5�5�5�5�5�5 6 6(646T6\6h6�6�6�6�6�6�6�6�67$7,787X7`7l7�7�7�7�7�7�7�7�7�7�78 8@8H8P8X8d8�8�8�8�8�8�8�8�8�89(909<9\9d9p9�9�9�9�9�9�9: :@:L:l:x:�:�:�:�:�:�:;$;,;8;X;`;h;p;|;�;�;�;�;�; < <,<L<X<|<�<�<�<�<�<�<�<�<�< ===4=@=`=l=�=�=�=�=�=�=�= > >(>4>T>\>h>�>�>�>�>�>�>�>�>?(?H?P?X?`?h?p?x?�?�?�?�?�?�? � �  000 0@0H0P0\0�0�0�0�0�0�0�0�0�0�0�011 1D1d1l1t1|1�1�1�1�1�1�1�1�1 2 2,2L2X2x2�2�2�2�2�2�233383D3d3p3�3�3�3�3�3�3�3 4444 4(40484D4d4p4�4�4�4�4�4�45 5@5H5T5t5|5�5�5�5�5�5 66,686X6d6�6�6�6�6�6�67747@7`7l7�7�7�7�7�7�7�78$8D8P8p8x8�8�8�8�8�8�89(949T9`9�9�9�9�9�9�9�9�9::(:H:P:X:d:�:�:�:�:�:�:�:;; ;,;L;X;x;�;�;�;�;�;�;�;<< <@<L<l<x<�<�<�<�<�<�<=(=H=T=t=|=�=�=�=�=�=�=�=>>$>D>L>X>x>�>�>�>�>�>�>�>�>�> ????$?D?P?p?|?�?�?�?�?�?�?   �   0(000<0\0h0�0�0�0�0�0�01181@1L1l1x1�1�1�1�1�1�1 2@2H2P2X2`2h2p2x2�2�2�2�2�2�2�2�2�2 3333<3H3h3t3�3�3�3�3�3484X4x4�4�4�4�4�4585X5x5�5�5�5�5 6 6@6`6�6�6�6�6�6�6777<7H7P7�7�7�7�7�7�7�7�7�7�7�7�7 8 8@8L8d8h8�8�8�8�8�8�89(949P9p9�9�9�9�9:,:0:L:P:p:�:�:�:�:�:   �    000$0<0d0h0�0�0�0�0101\1�1�1�1�12202P2p2t2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2343T3X3\3`3d3|3�3�3�3�3�3�3�3�3�3 444444444484<4X4x4�4�4�4�4�5�5�56@6\6�6�6�67<7p7�7�9�9�9�9:$:D:d:�:�:�:;0;h;�;�;<8<p<�<�<=8=\=t=�=�=�=>@>l>�>�>�>?<?l?�?�?�?     �   ,0\0�0�0�0�0�0101L1l1�1�1�1,2\2�2�2�2�2 3303`3�3�3�344h4�4�4 505\5�5�5�56P6�6�6�67<7p7�7�7�708h8�8�8�8�8 9L9P9T9p9�9�9:@:p:�:�:�: ; ;@;\;|;�;�; < <<<d<�<�<�<�<�<=4=X=t=�=�=�=>$>L>t>�>�>�>�> ?D?h?�?�?�?�?    �   0H0x0�0�0�001L1h1�1�1�1�1�1282X2x2�2�2�2 383X3p3�3�3�34D4d4�4�4�4�4 5$5H5l5�5�5�5�56(6D6d6�6�6�6�6�6747X7x=�=�=�=>,>`>�>�>�>?4?X?�?�?�?�?�?�?�?�?   (   000(0�0�0�0�0�0�0�0�0�0�0�0�0 111101`5X6`6d6�6�6�6�6�6�6�6�6�6�6l8t8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�89999j9n9r9v9|9�9�;�;�;�;�;�;�;�;�;<<
<<<<<<"<&<*<.<2<6<:<><B<F<J<N<R<V<Z<^<b<f<j<n<r<v<z<~<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<H=X=h=x=�=�=�=�=�=�=�=�=�=�>�> 0 �   p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1T2\2d2l2t2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23333$3,343z3~3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�5�5                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    