MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       "y��f��f��f�����g��A��~��A��	���e��f��0��A��&��A��g��A��g��Richf��                PE  L �ՐN        � !  �  �      ��     �                         P    z6                       � J   |� (     �                      @                                  � @            �                            .text   �s     �                   `.rdata  *0   �  @   �             @  @.data   �2   �      �             @  �.rsrc   �         �             @  @.reloc  p*      0                 @  B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �L$�A�	�Qf(��Y�f(��Y�f(��Y��X��X�W��Q�f.П��D�D$z�@� �@��x��^��Y��f(��YI�YA�H�@�������������̡$�V��H�QV�ҡ$��H�T$�AVR�Ѓ���^� ��̡$�V��H�QV�ҡ$��T$�H�D$�IRj�PV�у���^� �����������̡$��H�T$�I(��VWR�D$P�ы$��t$$���B�HV�ы$��B�HVW�ы$��B�P�L$Q�҃�_��^���̡$��P�D$���   ��P�D$$P�D$P�ҋL$�~ f��~@f�A�~@f�A����� �����̡$��Pd�D$P�D$PQ�J�у�� �̡$��Pd�D$P�D$P�D$PQ�Jt�у�� ������������̡$��PH�R,��`VW�D$P�ҋ��D$l�   ���_^��`� �̡$��P\�BXQ�Ѓ���������������̃�W��$��x�V�t$$�D$�L$�D$�P�RHW�D$P��h�  �����x��$��D$�D$W��D$�P�RH�D$Ph�  ���ҡ$��P�B0j h�  ������$��Q�B,���$h�  ���Ћ$��Q�B0jh�  ���Ћ$��Q�B0jh�  ������$��Q�B,���$h�  ���ЋL$$VQ���L  _^��� �������L  ����������̡$��P�B V�t$$����=mrict h'  ��Q  �$��Q��P�B8j���и   ^�  ������������QSVW���x �_xtKU3�9oh~B������D$t-�x uP��|  �D$���p�L$Q��|  �����ƉD$uӃ�;oh|�]S�|  3��wh�$��Bl�O �PQ�҉w ��W�`  ��_�F^[Y��̋D$V����  �WyN���F�$��zl+ƙ�����P�A �OP���D0 ��_^� �T$V��L$�D$P�FQ�NRP�h  ��t%�L$���T$�    t3��t�NPQ�N�yv  3�^� �;L$W�|$u�H��   _��    �V�NPR�Ev  �   ^� �����������̡$��I�PH���   Vj h�  Q�Ћ��D$�ȃ���  �yI���A+���������wq�$�� �T$���0Ɖ
�@�L$�^� �L$���T0Ɖ�P�D$�^� �T$���L0Ɖ
�@�L$�^� �L$���T0Ɖ��D$�^� �I k � � � ���̋D$�Ip�T$�@���R���\ �L��\H�T��\P�D$��f(��Y�f(��Y��X�f(��Y��X��%���Q�f/��v�D$f� f�Hf�P� �L$�!f/�v��L$�f/v�� W�f.���D�D${)�x��^��Y��Y��Y�� �H�P� �X�X�� ��������U������V��L$��  �M�Vj �D$PQ�NR�b  ��� �u�L$�2�  3�^��]� W��M�T$f(�f�f(�3���f�If�A~8�t$�*���X���Q�X��Q�Q��;��X��Q|��*�f.ȟ��D{I�x��^��	�Y��	�I�Y��I�I�Y��I�L$耣  �   ^��]� �A�A��L$�]�  �   ^��]� ̋T$V�r��u�D$��u�B+�^Ã��^�S�\$W3�3�3Ʌ�~�R;�����;΋�|���D$;�u�D$_[���^�_�C�[^���������������V�t$W�~��u�N�D$+�;�u_3�^�_��^�3�3�3҅�S�\$~�v;�����;׋�|���L$�T$���;�t�C[_^���������������V��������D$�L$PQ���G  ^� ���V�t$��蔻  ��u}�$����   ���   �҅��D$tF��tBjP���F�  �$����   �L$���   �Ѕ��L$u��@  3�^� ��@  �   @^� �$����   ���   �D$P�у�3�^� ������������U������dW�SVW���M�W�D$PQ�OR�D$,�D$$�D$�D$D�D$<�D$4�g  ��� �u3�_^[��]� �E�MW��4@�Gp����I���\0�L��\L0�D��\D0��f(��Y�f(��Y��X�f(��Y��X��Q�f.ߟ��Dz
f(�f(���%x��^�f(��Y��Y��YċGp�M�I�,��\,0�\��\\0�d��\d0��f(��Y�f(��Y��X�f(��Y��X��Q�W�f.���Dzf(�f(��T$@�&�x��^�f(��Y��t$@�Y��Y�f(��T$f(��Yd$ �YL$f(��YD$�Y��\��l$ �Y��\��D$`f(��Y��|$ �\�f(��Y�f(��Y��YT$@�\��L$@�Y��|$�Y��\��X�f(��X��Y��\��XL$`f(��Y�f(��Y��X�f(��Y��X�W��Q�f.ܟ��Dzf(�f(�f(���%x��^�f(��Y��Y��YӋ]�M�D$(Pf�Qf�K��f�S������������p�L7�\L$0�[�7�\D$(�#�T7�k�\T$8�f(��Y�f(��Y�f(��Y��X��X�W�f/�v*���f(�f(��\�f��\��\�f�Sf�C_^�   [��]� �������SV�t$�V3���W~�>�\$��9t����;�|�_^3�[�PV��������L$ ��_^��   [���������SV�t$�V3���W~�>�\$��9t����;�|�_^3�[�PV�������L$ ��_^��   [���������V������"����N�*�  ��^�"@  �̡$��H�A��  SUV�T$WR�Ћ$��Q�J3�Wj��D$h(�P�эT$$R�� �$��H�A�T$(R�Ћ$��Q��$�  �B`��W���Ћ�����o��  ���$��Q�BtV���Ћ$�W�|$4�|$<���   �JP�D$8P�ы$����   �P�L$<Q�҃�=   ��  ��  =�   �!  ���1 �$�H1 Wh���$(  �
���Wh���$h  �������$   Q��$�  VR�"���P��$p  P��$�  Q�;  ��P��$�  R�;  P�� �$��H�A��$   R�Ћ$��Q�J��$�  P�ы$��B�P��$  Q�ҡ$��H�A��$|  R�Ћ$��Q�J��$@  P�у�$�8  Wh���$H  �/���Wh���$�  ������$@  R��$T  VP�G���P��$�  Q��$$  R��:  ��P��$X  P�:  P�� �$��Q�J��$`  P�ы$��B�P��$$  Q�ҡ$��H�A��$h  R�Ћ$��Q�J��$�  P�ы$��B�P��$`  Q�҃�$�\  Wh����$h  �S���Wh���$  �A�����$`  P��$T  VQ�k���P��$  R��$�  P��9  ��P��$8  Q��9  P� �$��B�P��$@  Q�ҡ$��H�A��$�  R�Ћ$��Q�J��$h  P�ы$��B�P��$  Q�ҡ$��H�A��$�  R�Ѓ�$�  Wh���$�  �x���Wh���$  �f�����$�  Q��$�  VR����P��$  P��$�  Q�
9  ��P��$  R��8  P�3 �$��H�A��$   R�Ћ$��Q�J��$�  P�ы$��B�P��$�  Q�ҡ$��H�A��$  R�Ћ$��Q�J��$�  P�у�$�  Wh���$�  ����Wh���$(  ������$�  R��$�  VP����P��$0  Q��$�  R�/8  ��P��$�  P�8  P�X �$��Q�J��$�  P�ы$��B�P��$�  Q�ҡ$��H�A��$�  R�Ћ$��Q�J��$<  P�ы$��B�P��$�  Q�҃�$��  WhԒ��$�  �����Wh���$�  ������$�  P��$4  VQ�����P��$�  R��$�  P�S7  ��P��$�  Q�B7  P�| �$��B�P��$�  Q�ҡ$��H�A��$�  R�Ћ$��Q�J��$H  P�ы$��B�P��$�  Q�ҡ$��H�A��$�  R�Ѓ�$��  WhĒ��$�  �����Wh���$H  �������$�  Q��$  VR�����P��$P  P��$�  Q�x6  ��P��$�  R�g6  P� �$��H�A��$   R�Ћ$��Q�J��$�  P�ы$��B�P��$(  Q�ҡ$��H�A��$\  R�Ћ$��Q�J��$   P�у�$�  Wh����$8  ����Wh���$  �������$0  R��$�  VP�#���P��$   Q��$D  R�5  ��P��$x  P�5  P�� �$��Q�J��$�  P�ы$��B�P��$D  Q�ҡ$��H�A��$�  R�Ћ$��Q�J��$,  P�ы$��B�P��$P  Q�҃�$�8  Wh����$x  �/���Wh���$X  ������$p  P��$$  VQ�G���P��$`  R��$  P��4  ��P��$�  Q�4  P��
 �$��B�P��$�  Q�ҡ$��H�A��$  R�Ћ$��Q�J��$8  P�ы$��B�P��$l  Q�ҡ$��H�A��$�  R�Ѓ�$�]
  Wh����$�  �T���Wh����$�  �B���Wh���$�  �0����$����   �JH�D$0P�у���$�  RP��$�  P��$�  VQ�8���P��$�  R��$�  P�3  ��P��$�  Q�3  ��P��$l  R�3  ��P��$H  P�3  P�	 �$��Q�J��$P  P�ы$��B�P��$t  Q�ҡ$��H�A��$�  R�Ћ$��Q�J��$�  P�ы$��B�P��$�  Q�ҡ$��H�A��$�  R�Ћ$��Q�J��$�  P�ы$��B�P��$�  Q�҃�0��  Wh����$8  �����Wh����$  �����Wh���$�  �����$����   �AL�T$0R�Ѓ���$0  Q��$�  R����  P��$  P��$l  VQ����P��$  R��$\  P�12  ��P��$0  Q� 2  ��P��$  R�2  ��P��$�  P��1  P�8 �$��Q�J��$�  P�ы$��B�P��$  Q�ҡ$��H�A��$8  R�Ћ$��Q�J��$\  P�ы$��B�P��$�  Q�ҡ$��H�A��$�  R�Ћ$��Q�J��$  P�ы$��B�P��$<  Q�ҡ$��H�A��$`  R�Ѓ�4�T  Whp���$x  �K���Wh���$X  �9�����$p  Q��$�  VR�c���P��$`  P��$�  Q��0  ��P��$�  R��0  P� �$��H�A��$�  R�Ћ$��Q�J��$�  P�ы$��B�P��$�  Q�ҡ$��H�A��$l  R�Ћ$��Q�J��$�  P�у�$�y  Wh`���$�  �p���Wh���$�  �^�����$�  R��$D  VP����P��$�  Q��$4  R�0  ��P��$  P��/  P�+ �$��Q�J��$  P�ы$��B�P��$4  Q�ҡ$��H�A��$X  R�Ћ$��Q�J��$�  P�ы$��B�P��$�  Q�҃�$�  �$��H�A��$�   R�Ћ$��Q�JWj���$�   hP�P�ы$��B�P��$  Q�ҡ$��H�AWj���$  h�R�Ћ$��Q�J(��$�  VP�ы$����B�P��$�   Q�ҡ$��H�A��$�   RV�Ћ$��Q�J��$�  P�ы$��B�P��$�   ��@Q�ҡ$��H�I�T$dR��$�   P�ы$��B�P<���L$`�ҋ$��Qj��RLj���$�   QP�L$p�ҡ$��H�A��$�   R�Ћ$��Q�R��$�   P�L$hQ�ҡ$��P�B<����$�   �Ћ$��Q�RLj�j���$�   QP��$�   �ҍ�$�   P� �$��Q�J��$�   P�ы$��B�P�L$hQ�ҡ$��H�A��$�   R�Ћ$��Q�J��$   P�э�$�   �  =  ��  =@B ��  �$��H�A��$�   R�Ћ$��Q�JWj���$�   h8�P�ы$��B�P��$�   Q�ҡ$��H�AWj���$�   h�R�Ѝ�$�  VQ�^����$����B�P��$�   Q�ҡ$��H�I��$�   R��$�   P�ы$��B�P<��<�L$p�ҋ$��Qj�j�VP�BL��$�   �Ћ$��Q�J�D$@P�ы$��B�@�L$DQ�T$xR�Ћ$��Q���B<�L$@�Ћ$��Q�RLj�j���$�   QP�L$P�ҍD$@P�` �$��Q�J�D$DP�ы$��B�P�L$xQ�ҡ$��H�A��$�  R�Ћ$��Q�J��$�   P�э�$�   ��  �$��H�A�T$ R�Ћ$��Q�JWj��D$,h$�P�ы$��B�P��$�   Q�ҡ$��H�AWj���$�   h�R�Ћ$��Q�J(��$�  VP�ы$����B�P��$�   Q�ҡ$��H�A��$�   RV�Ћ$��Q�J��$�  P�ы$��B�P�L$P��@Q�ҡ$��H�I�T$R��$�   P�ы$��B�P<���L$�ҋ$��Qj��RLj���$�   QP�L$ �ҡ$��H�A�T$PR�Ћ$��Q�R�D$TP�L$Q�ҡ$��P�B<���L$P�Ћ$��Q�RLj�j��L$(QP�L$`�ҍD$PP�  �$��Q�J�D$TP�ы$��B�P�L$Q�ҡ$��H�A��$�   R�Ћ$��Q�J��$�   P�эL$4�$��B�PQ�҃��$����   ��T$0R�Ћ$��Q�B`��U���Ћ�������C����$��Q�J�D$ P�ы$��B�PWj��L$,h�Q�ҍD$4P��  �$��Q�J�D$8P�у�_^][�Ġ  Ë��  [  6! " �" �# �$ % Z& �' c) >* �0  	
���������̃�V��L$�r  �L$ �Vj �D$PQ�NR�iG  ��� ��L$tO�t$�D$ PVQ��������� �t&�D$ ;D$u7�T$$R�D$VP���������� �u!�L$�q  �L$�Ȉ  3�^��� �L$$��L$�q  �L$览  �   ^��� ����������̋T$�D$ SU�l$VW�|$ �ٍL$ QWUR���    �����t$ ;t$�D$$�L$,�0�9t@�D$,�T$RPWVU���k����|$ t1�L$,�9�T$ RWUV��������t$ ;t$t(;t$u�_^]�   [�  �D$0_^]�     �   [�  _^]3�[�  ����U������|SVW��3ۉ_h�_x�$����   ���   ��;ÉD$u&�$����   ���   �T$R�Ѓ�3�_^[��]� �OtjP讑  �$����   �L$���   �Ѕ�u*�$����   ���   �D$P�у��   _^[��]� �$����   �L$���   S�ҋȉG��  �ȉG�K ���g  �G�$��Q\P�BX�ЉGl�G�$��QHh�  P���   �ЉGh�G�$��QHSh�  P���   �ЉGp�G�$��QHh�  P���   �Ћ$��QH���GSh�  P���   �ЋW�R��,SV�OP�GhP�҅�u�L$�Z%  3�_^[��]� �?  ;ÉGt��OSQ���G@  ��tЋOh�$��B���   hP���h�  Q�҃�;ÉGxt��D$HP�L$dQ�O3�S�1 ����  ���$    �t$`��;t$H�\$$�t$\��  ��$    V���������m  �T$XR�D$hPV���^����$��Q���   hP�h  h�   �Ћ����������$��Q���   hP�h  h�   �Ћ؃��ۉ\$T������$��Q���   hP�h  j(�Ѓ���������L$d�T$X��P��F ��C�Gx�<� ��u7�0�_p�I�~ÍËGx����f� �~Cf�@�~C�\$Tf�@�� �@�p�Gx���p�Gx���A�Ox�<� ��u3��Op�R�~����Gx����f� �~Af�@�~Af�@���A�X�Ox���t$\�X�Ox���B��;t$H�t$\�r����\$$�O�T$HR�D$dPS�[ ���3����h �D$$    ��   ��Ox�T$$������   �{ ��   �3�Ox����J���N�Wx�N���R���~�Vu�Wx��92u�R��V�~u�Wx��92u�R��V�T$dRQ�OP�GP�lE  �L$d��t���������N�P�V�F$    ��F$   ��N�W�OPR�-S  �[���D����D$$��;Gh�D$$�����h �H�Wҍ_8�OH�\$D��L$8��W@�WP�D$$    ��  ��Ox�T$$�<� ����  � ��{ ��  �{��  �S��L$hQ�ORPQ�O�\$|�D  �L$h��t���#����q�H�L$\�
3��D$\������OP�GP�T$`�t$l�IR  �T$\�L$X�%���T$(2��D$   �t$ �T$�I �4������D$0�Gx�t$�4�3��{ �D$,�D$4��  ���D$���C u'9D$ u!9C$�K�D$   uN�C�D$(�D$    �=�{$ u7��t�|$  u,�C;�u�C�D$(�D$    ��K9L$(u�K�D$   �|��F  �\��T$9����D$<�D$@3�9D$�T$�D$P�D$T��   �T$PR�T$@R�T$pR���T$8R�T$(Q�L$D�D$`� PQR��������������D$,�L$L;tD���   R�T$�O@Q�L$LQRP��$�   P���v����~ f�F0�~@f�F8�~@f�F@�#�T$<�N0Q�L$RP�D$<PQ����������A����%���|$  ��   �T$���L$TQ�T$DR�L$pQ�L$4�T$@R�Q�L$,�D$`�D$DRPQ���������������D$4�T$L;tD�T$8���   Q�OPQ�L$ RQP��$�   R�������~ f�FH�~@f�FP�~@f�FX�#�T$@�NHQ�L$RP�D$<PQ���5������z����%���|$ ��   �{$ ��   �|$T ��   �C9D$@u�C�L$�T$,R��P�D$ PR���>������#����L$D�T$���   P�G@P�D$4QRP��$�   Q��������~ �%��f�F0�~@f�F8�~@f�F@�  ݆�   f(��\FHf(��\NPf(��\VXݞ�   f�F0f�N8f�V@��   �|$  ��   �{$ ��   �|$P t�C9D$<u�C�L$�T$4R��P�D$ PR���e������J����L$8�T$���   P�GPP�D$<QRP��$�   Q�������~ �%��f�FH�~@f�FP�~@f�FX�6݆�   f(��\F0f(��\N8f(��\V@ݞ�   f�FHf�NPf�VX�V8�^@���   �T$@�D$P�Y��YًL$<f(��YF0�XF�N �X��V(f�F`f�Nh���   �X�f�Vp�FH�VP�^X�T$(�T$T�Y��Y��XF�Y��N �D$�X��V(f�Fxf֎�   �T$ �T$���X�f֖�   �4������D$0�Gx�t$�4�3��{ �D$,�D$4�A�����  �|$ �\$te�D$0�T$,RQSP���������������T$D���   Q�G@P�D$4RSP��$�   Q�������~ �%��f�F0�~@f�F8�~@f�F@�|$  ti�D$(�L$0�T$4RPSQ���^������C����L$4���   R�GPP�D$@PSQ��$�   R�������~ �%��f�FH�~@f�FP�~@f�FX�|$ u8݆�   f(��\FHf(��\NPf(��\VXݞ�   f�F0f�N8f�V@�=�|$  u6݆�   f(��\F0f(��\N8f(��\V@ݞ�   f�FHf�NPf�VX�F0�V8�^@���   �Y��Y��XF�Y��N �X��V(f�F`���   f�Nh�X�f�Vp�NH�VP�^X�Y��Y��Y��F�X��N �X��V(f�Fx�X�f֎�   f֖�   �D$\�\$l�L$X�D$(�D$d�D$ �D$��<�C  �D$   �D$�����W��H��D$$��;Gh�D$$�����\$D�L$8�	�@�f.ȟ��Dz�f.ȟ��D�	z����#f.����Dz��GPf.��Dz �G@f.��D�GPz �_@�_P��O@f.ʟ��Dz�G@3�9wh��   �I �Ox�<� t{�$��B�M���   j h�  �҅�t8�Gx�����   �^G@���   �Ox�����   �^GP���   �$�Wx���x����   �Ox�����   ��;wh�p�����p��D$8�Y����Y���$����   ���   �T$R�Ѓ�_^�   [��]� ���U������xVW�������EP���s����L$l�� W��}�F0�F   �$��Q���   j hxvpi���Ћ$��Q�*����   j hyvpi���D$`�Ћ$��Q�}�*����   j h�  ���D$X����$��Q���$�D$<���   h�  �����\$8�$���Q���   ���$h�  �����T$@�������v����D$@���f/D$8v�D$8�D$P�Mj���\$�D$l�$h �  �VW  �L$lQ�M�T$dR�D$PP�W  ���*  �D$H�Y���YD$@�XF0�F0�$��Q���   j haqpi�L$t�Ћ$��Q�����   j haqpi�L$t���к   #��  ���  �F03�f/���~$��   9Nh��  �d$8�Vx�<� ����   �|$4 � ���   �YF0���   t8�Fx������   ���   �\�f/�r�����   �\����   �Vx�����   �P8�X@�Y�f(��YH0�Y��@�X��H �X��P(�Fp�f� �X�f�Hf�P����;Nh�4������+  9Nh��   �d$8�5���-p�3��Fx�<� ����   �|$4 � ���   �YF0f(��\����   t=�Vx�����   ���   ��fT��\�f/�r�����   �\����   �Fx�����   �PP�XX�Y�f(��YHH�Y��@�X��H �X��P(�Fp�f� �X�f�Hf�P����;Nh�'������*  ���W  �F0f/��r�   �3�9V$t��3��~(�V$�$��B�V(�@,3ыM���*��$h�  ��3�9N(t~9Nh��  3ҍI �Fx�<� ��tT� ���   �YF0�H0�P8�X@�Y��Y��XH�Y��@ �X��P(�Fp�f��X�f�@f�P����;Nh|��k  9Nh�b  3���I �Fx�<� ��tX� ���   �YF0�HH�PP�XX�Y��Y��Y��@�\��H �\��P(�Fp�f� �\�f�Hf�P����;Nh|���  W�3�f/F0�F$   ��   9Nh��  �-���%p�3��Vx�<� ����   �|$4 � ���   �YF0���   t4�Fx������   fT�f/��   r��f(��\��   ���   �Vx�����   �P8�X@�Y�f(��Y@0�X@�Y��H �X��P(�Fp�f� �X�f�Hf�P����;Nh�<�����   9Nh��   3���    �Fx�<� ����   �|$4 � ���   �YF0���   t)�Vx�����   f/��   ��r��݂�   ݚ�   �Fx�����   �HH�PP�XX�Y��Y��Y��@�\��H �\��P(�Fp�f� �\�f�Hf�P����;Nh�C�����$��Q�M�B,���$h�  �Ћ$����   �N�Bj j���F0�$��Q�M�B,���$h�  ��j j j hed�����  j h�  ���  ���L$lQ�M�T$dR�D$PP�XQ  ��������}�M�tQ  ��t
�Ntj �%�  j �F    �g�  ��������W�W���F0������L$l� _�   ^��]� �������VW��������|$�GP�������Gt�NQ�j(�u�  ��� �u_^� �$���B�O���   ���$h�  ���^0�$��P�O���   j h�  ��3Ʌ��   �F0f/����   9Nh�
  3Ґ�Fx�<� ��tP� �F0�P8�X@�Y�f(��YH0�Y��@�X��H �X��P(�Fp�f� �X�f�Hf�P����;Nh|�j �"�  ��_�   ^� 9Nh��  3ҋFx�<� ��tP� �F0�HH�PP�XX�Y��Y��Y��@�\��H �\��P(�Fp�f� �\�f�Hf�P����;Nh|�j ��  ��_�   ^� W�f/F0��   9Nh��   3ҍ�    �Fx�<� ��tL� �N0�@0�P8�X@�Y��Y��X@�Y��H �X��P(�Fp�f� �X�f�Hf�P����;Nh|�j ��  ��_�   ^� 9Nh~k3ҋ��Fx�<� ��tP� �F0�HH�PP�XX�Y��Y��Y��@�\��H �\��P(�Fp�f� �\�f�Hf�P����;Nh|�j ��  ��_�   ^� �����U������SVW�������EP��������}���x�  �NQj(��諌  ��脌  3�9Nh�]  �]���3ҋFx�<� �<��1  ���  ����   �Hx�\H`���   �\Ph���   �\Xpf(��Y�f(��Y��X�f(��Y��X��Q�f(�f.5�����Df(��Y%��{�-x��^��Y��Y��Y݋�Y��Ỹ�`�Y�� �X��H�X��P�XӋFp�f� f�Hf�P�a  ���   ���   ��X��Y��f/��  ���   ��-�  �\���   ����   ���  �Y���Fx���p8�x@f(��Yh0�Y��Y�f(��\PH�Y�f(��\XP�Y�f(��\`X�Y��H�X��P �X��X(�X��X��X��X��  �Fx��f(��\PHf(��\XPf(��\`X�2  �Fx���X8�`@�Y�f(��YP0�XP�Y��H �X��X(�Fp�f��X�f�H�  ���   ��-�  �\���   ����   ����   �Y���Fx���hH�pP�xXf(��\P0�Y��XPf(��\`@�Y��Y��Y��d$ f(��P(�XT$ �Y�f(��\X8�Y��H �X��X��X��X�������Fx��f(��\P0f(��\X8f(��\`@��Fx���PH�XP�`X�Y��Y��Y��H�X��P �X��X(�X܋Fp�f�f�Pf�X����;Nh������$����   �N�Bj j��j ��  j h�  ���  ��_^[��]� �����V�t$��W��u_3�^� ���&�  ��uhShҝ V�wt�rI  �؃���tH��肈  �GPj(��赈  ��莈  �L$ �T$�D$QRPS��������t[_�   ^� �������[_3�^� _�   ^� ��������������̃�VWhP�h�  hp�h�   �C  ������t���  �N����t�  �3��$��H�A�T$R�Ћ$��Q�Jj j��D$h��P�у��T$R�L$��  �8Vh'  ��  ��PWh(  h'  ��  ��Phҝ �J  ���L$���t�  �$��H�A�T$R�Ѓ�_��^���������̋D$S�\$VW�|$PWS���  3�;�� �u_^3�[� �N�N(�Nx�Nh�NW�Ή^t�J���_^�   [� ���������������S�\$��V�t$W��u=j ���5 � G�����w(j ���  � �L$�T$PQR�������_^�   [� �D$�L$VSPQ���NG  _^[� �����������������������U�����E��l  �SVW��t:�u6�$����   ���   �҅��D$u&�$����   ���   �T$R�Ѓ�3�_^[��]� �MjP�Xr  �$����   �L$���   �Ѕ�u�L$�  �   _^[��]� �$����   �L$���   j �ЋN;��}u�̑  ��蕾��9Flt������W��������N0W�f/��x�v�NX�F`�
�N`�FX�~ u#�$��Q���   j h�  ��������؉F$��$   j/Q���  �x����T$Rh�  �D$0P���D$,�D$$�D$�����x��L$Qh�  �T$HR���D$,�D$$�D$�����N��$  P�z����$��Qd�}�JpP�FPW�ы$��L$Q�D$    �D$(   �Bd���   h�  W�ҡ$����   ��T$(R��3ۃ�9^h��  �Nx�<� ��  �$��Bd�H`jW�ыF$���� j �#  ���   �~( ����   �T$,R�w����Fx�NX����P8�X@�Y�f(��Y@0�X@�Y��H �X��P(�X��D$�L$�T$ �j �T$R��P���2���j �L$DQ�������Vx���H0�P8�X@�F`���Y��Y��Y��@ �\��P(�\��X�\���$�   ��$�   ��$�   �	j ��$�   ��PQ��讻���Y  �T$DR�����Fx�F`����PP�XX�Y��Y�f(��@ �YHH�X��P(�X��X�X���$�   ��$�   ��$�   �j ��$�   R��P���*���j �L$,Q��������Vx���HH�PP�XX�FX���Y��Y��Y��@ �\��P(�\��X�\��\$X�D$`�T$h�	j �D$\��PQ��貺���]  �$��Bd�P�L$DQW�ҋFx�F`�$�����H0�P8�X@�Y��Y��Y��@ �\��P(�\��X��$�   ��$  �\���$�   �Bd�	j ��$�   R�Pt��QW�ҡ$��Hd�Aj �T$HRW�ЋNx���PP�XX�FX�$����Y��Y�f(��@ �YHH�\��P(�\��X�\���$�   ��$�   ��$�   �Bd��$�   �1  �$��Hd�A�T$,RW�ЋNx�����   �H0�P8�X@�YFX�X��   �$����Y��Y��XH�Y��@ �X��P(��$�   ��$�   �X���$�   �Bd�	j ��$�   R�Pt��QW�ҡ$��Hd�Aj �T$`RW�ЋNx�����   �HH�PP�XX�YF`�X��   �$����Y��Y��Y��@ �X��P(�X��X�X���$�   ��$�   ��$�   �Bd��$�   �	j R�Pt��QW�҃�8�$��Hd�Aj ��$  RW�Ћ$��Qd�B`jW�Ћ$��Qd�Fx�����   j j��QW�҃�$��;^h�����$��Hd�Q`j W�ҡ$��T$R�D$   �D$$   �Hd���   h�  W�Ћ$����   �
�D$$P�ы$����   ���   �L$$Q�҃�_^�   [��]� �������������̡$�V�񋈈   ���   V�҃��    ^��������������̡$��H�QV�t$V�ҡ$��H�T$�AVR�Ћ$��Q�B<�����Ћ$��Q�L$�RLj�j�QP���ҋ�^���������̸ҝ ����������̡$��H�QV�t$V�ҡ$��H�Qj j�h��V�҃���^� �������������V������r����N�z�  ���s  �D$t	V�8  ����^� ������������̃�������u��á$��H�A�$R�Ћ$��Q�Jj j��D$hd�P�эT$R�	�  �$��H�A�T$R�Ћ$��Q�J�D$P�ы$��B�Pj j��L$(h(�Q�ҍD$0P��  �$��Q�J�D$4P�ы$��B�P�L$8Q�ҡ$��H�Aj j��T$Dh�R�ЍL$L��LQ�p�  �$��B�P�L$Q�ҡ$��H�A�T$R�Ћ$��Q�Jj j��D$h��P�эT$R�%�  �$��H�A�T$ R�Ћ$��Q�J�D$$P�ы$��B�Pj j��L$0h(�Q�ҍD$8P���  �$��Q�J�D$<P�ы$��B�P�L$@��@Q�ҡ$��H�Aj j��T$hd�R�ЍL$Q��  �$��B�P�L$Q�҃��   �������������������������������̋D$�� t��t3�ù(���  �����ø   ���������U��E�$�� ]�̋�� l����������l����������̅�t��j�����̡$��P��  ��$��P��(  ��U��$��P��   ��V�E�P�ҋuP��説  �M���  ��^��]� ��������̡$��P��$  ��U��$��H��  ]��������������U��$��H���  ]�������������̡$��H��  ��U��$��H���  ]��������������U��$��H��x  ]��������������U��$��H��|  ]��������������U���EV���l�t	V��4  ����^]� ��������������U��$��PH�EPQ���  �у�]� �U��$��P�B4VW�}j��h�  ���ЋMWQ����8  _^]� ��������������U��V���PXW�ҋ}P�����  ���Et�_�   ^]� �M�UPWQR����9  _^]� �����������U��S�]VW��j ����  �8�  �}uI�~ uC�$��P���   j h�  ���Ѕ�u�$��QP���   h�  ���Ѕ�t	_^3�[]� �M�U�EQ�MRPSWQ���_9  _^[]� ��������U��EP�A    ��  ��]� �����̸   �A� ������A   � ������U���@S�]��`��VW��u�G   �}  ����   �M3�V��  �8�  u4��v  P�w�T  �$��P�M�B4��jh�  ��_^�C�[��]� �MV�e�  �8�  u�E�M��RPQ����_^�   [��]� �MV�5�  �8�  t�MV�$�  �8��  �$��P�M�B4jh�  �Љw�  ����  �E�H��BXj	��P����3��؃�;މu�t�$��QH���  VS�Ѓ��E��M�;O�f  9w�]  �$��B�M���   Vh�  �҅�u!�$��P�M���   Vh�  �Ѕ��  �$��Q�M�B4Vh�  ��;�t
V���������E��G�$����   ���   �Ћ];މE���   ;���   S��|  �M���jQ�ˉu��uĉuȉủuЉu؉u��b  �U�E��ˉu��u�u�U�E��]��E�   ��q  ��t!��t��t�u���E�   ��E�   ��E�   �Z�  �M�;�t�v  ��BX�M�Q����P�+�  �M܃�;�t�v  �M��t�  �M��l�  �M������]�M�U�EQSRP���6  _^[��]� �M������_^�   [��]� ��������������U��$��P�E���   ��VWP�EP�E�P�ҋu���$��H�QV�ҡ$��H�QVW�ҡ$��H�A�U�R�Ѓ�_��^��]� ������������U��E��u�(��MP�EPQ��  ��]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3hp�j;hp�j�]0  ����t
W���^�  �3����Fu_^]� �~ t3�9_��^]� �$��H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   �$��H<�Q��3Ʌ����^��������������̃y t�   ËA��uË$��R<P��JP�у��������U����u�$��H�]� �$��J<�URP�A�Ѓ�]� ���������������U��(���u�$��H�]Ë$��J<�URP�A�Ѓ�]�U��(���$��Vu�$��H�1��$��J<�URP�A�Ѓ����$��Q�J�E�SP�ы$��B�P�M�QV�ҡ$��H�A�U�R�Ћ$��Q�Jj j��E�h��P�ы$��B�@@�� j �M�Q�U�R�M��Ћ$��Q�J���E�P���у���[t.�$��B�u�HV�ы$��B�P�M�Q�҃���^��]á$��P�E��RHjP�M��ҡ$��P�E�M��RLj�j�PQ�M��ҡ$��H�u�QV�ҡ$��H�A�U�VR�Ћ$��Q�J�E�P�у���^��]���������������U��(���$��SVu�$��H�1��$��J<�URP�A�Ѓ����$��Q�J�E�P�ы$��B�P�M�QV�ҡ$��H�A�U�R�Ћ$��Q�Jj j��E�h��P�ы$��B�@@�� j �M�Q�U�R�M��Ћ$��Q�J���E�P���у���t/�$��B�u�HV�ы$��B�P�M�Q�҃���^[��]á$��P�E��RHjP�M��ҡ$��P�E�M��RLj�j�PQ�M��ҡ$��H�A�U�R�Ћ$��Q�Jj j��E�h��P�ы$��B�@@��j �M�Q�U�R�M��Ћ$��Q�J���E�P���у����3����$��P�E��RHjP�M��ҡ$��P�E�M��RLj�j�PQ�M��ҡ$��H�u�QV�ҡ$��H�A�U�VR�Ћ$��Q�J�E�P�у���^[��]����������������U��(���$��SVu�$��H�1��$��J<�URP�A�Ѓ����$��Q�J�E�P�ы$��B�P�M�QV�ҡ$��H�A�U�R�Ћ$��Q�Jj j��E�h��P�ы$��B�@@�� j �M�Q�U�R�M��Ћ$��Q�J���E�P���у���t/�$��B�u�HV�ы$��B�P�M�Q�҃���^[��]á$��P�E��RHjP�M��ҡ$��P�E�M��RLj�j�PQ�M��ҡ$��H�A�U�R�Ћ$��Q�Jj j��E�h��P�ы$��B�@@��j �M�Q�U�R�M��Ћ$��Q�J���E�P���у����3����$��P�E��RHjP�M��ҡ$��P�E�M��RLj�j�PQ�M��ҡ$��H�A�U�R�Ћ$��Q�Jj j��E�h��P�ы$��B�@@��j �M�Q�U�R�M��Ћ$��Q�J���E�P���у���������$��P�E��RHjP�M��ҡ$��P�E�M��RLj�j�PQ�M��ҋu�E�P�������$��Q�J�E�P�у���^[��]�������U��(���$��SVu�$��H�1��$��J<�URP�A�Ѓ����$��Q�J�E�P�ы$��B�P�M�QV�ҡ$��H�A�U�R�Ћ$��Q�Jj j��E�h��P�ы$��B�@@�� j �M�Q�U�R�M��Ћ$��Q�J���E�P���у���t/�$��B�u�HV�ы$��B�P�M�Q�҃���^[��]á$��P�E��RHjP�M��ҡ$��P�E�M��RLj�j�PQ�M��ҡ$��H�A�U�R�Ћ$��Q�Jj j��E�h��P�ы$��B�@@��j �M�Q�U�R�M��Ћ$��Q�J���E�P���у����3����$��P�E��RHjP�M��ҡ$��P�E�M��RLj�j�PQ�M��ҡ$��H�A�U�R�Ћ$��Q�Jj j��E�h��P�ы$��B�@@��j �M�Q�U�R�M��Ћ$��Q�J���E�P���у���������$��P�E��RHjP�M��ҡ$��P�E�M��RLj�j�PQ�M���j h���M�袢���$��P�R@j �E�P�M�Q�M��҅��$��H�A�U�R���Ѓ���t/�$��Q�u�BV�Ћ$��Q�J�E�P�у���^[��]Ë$��M��B�PHjQ�M��ҡ$��P�E�M��RLj�j�PQ�M��ҋu�E�P���ˡ���$��Q�J�E�P�у���^[��]���������������U��$��H<�A]����������������̡$��H<�Q�����V��~ u>���t�$��Q<P�B�Ѓ��    W�~��t���ʛ  W�$  ���F    _^��������U���V�E�P���ޮ  ��P��������M��艛  ��^��]��̃=0� uK�(���t�$��Q<P�B�Ѓ��(�    �4���tV���@�  V�*$  ���4�    ^������������U���8�$��H�AS�U�V3�R�]��Ћ$��Q�JSj��E�h��P�ы$��B<�P�M�Q�ҋ�$��H�A�U�R�Ѓ�;�u^3�[��]�V�M�]���  �M�Q�U�R�M��X�  ����   W�}�}���   �$����   �U��ATR�Ћ�����tB�$��Q�J�E�P���у��U�Rj�E�P�������$��Q�ȋBxW�Ѕ��E�t�E� ��t�$��Q�J�E�P����у���t�$��B�P�M�Q����҃��}� u"�E�P�M�Q�M���  ���;����E�_^[��]ËU��U�_�E�^[��]��������������U���DSV�u3�;�]�u_�$��H�A�U�R�Ћ$��Q�JSj��E�h��P�ы$��B<�P�M�Q�ҋ�$��H�A�U�R�Ѓ�;�u^3�[��]�V�M�]���  �M�Q�U�R�M����  ���p  W�}��I �E����   �$����   �U��ATR�Ћ�������   �$��Q�J�E�P���ы$��B���   ���M�Qj�U�R���Ћ$��Q�J���E�P�ы$��B�P�M�QV�ҡ$��H�A�U�R�Ћ$��Q�Bx��W�M��Ѕ��Et�E ��t�$��Q�J�E�P����у���t�$��B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*�$����   P�BH�Ћ$��Q���ȋBxW�Ѕ�t"�M�Q�U�R�M��r�  ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M����  �EP�M�Q�M�u��u��  ����   �u���E���tA��t<��uZ�$����   �M�PHQ�ҋ$��Q���ȋBxV�Ѕ�u-�   ^��]Ë$����   �E�JTP��VP�[�������uӍUR�E�P�M���  ��u�3�^��]����������V��~ u>���t�$��Q<P�B�Ѓ��    W�~��t��芖  W�t  ���F    _^��������h8�Ph� ��  ���������������h8�jh� ��  ����uË@����U��V�u�> t/h8�jh� �S�  ����t��U�M�@R�Ѓ��    ^]���U��Vh8�jh� ����  ����t�@��t�M�UQR����^]� 3�^]� ���U��Vh8�jh� �����  ����t�@��t�M�UQR����^]� 3�^]� ���U��Vh8�jh� ����  ����t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������Vh8�jh� ���L�  ����t�@��t��^��^��������U��Vh8�j h� ����  ����t�@ ��t�MQ����^]� ��������������U��Vh8�j$h� �����  ����t�@$��t�M�UQR����^]� 3�^]� ���U��Vh8�j(h� ����  ����t�@(��t�M�UQR����^]� 3�^]� ���U��Vh8�j,h� ���Y�  ����t�@,��t�M�UQR����^]� 3�^]� ���U��Vh8�j0h� ����  ����t�@0��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh8�j4h� �����  ����t �@4��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh8�j8h� ���y�  ����t%�@8��t�M�E�UQ�M���$RQ����^]� 3�^]� ������U��Vh8�j@h� ���)�  ����t�@@��t�M�UQR����^]� 3�^]� ���U��Vh8�jDh� �����  ����t�@D��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh8�jHh� ����  ����t �@H��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh8�jLh� ���I�  ����t�@L��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh8�jPh� �����  ����t�@P��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh8�jTh� ����  ����t �@T��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh8�jXh� ���Y�  ����t �@X��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh8�jdh� ���	�  ����t%�@d��t�E�M�U���$Q�MRQ����^]� 3�^]� ������U��Vh8�jhh� ����  ����t �@h��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh8�jlh� ���i�  ����t$�@l��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh8�jph� ����  ����t �@p��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh8�jth� �����  ����t�@t��t�M�UQR����^]� 3�^]� ���U��Vh8�jxh� ����  ����t �@x��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh8�j|h� ���9�  ����t�@|��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh8�h�   h� �����  ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh8�h�   h� ����  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh8�h�   h� ���F�  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh8�h�   h� �����  ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh8�h�   h� ����  ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh8�h�   h� ���V�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h�   h� ����  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h�   h� ����  ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh8�h�   h� ���f�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h�   h� ����  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h�   h� �����  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h�   h� ���v�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h�   h� ���&�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h�   h� �����  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh8�h�   h� ����  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh8�j\h� ���9�  ����t�@\��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh8�j`h� �����  ����t�@`��t�M�UQR����^]� 3�^]� ���U��Vh8�j<h� ����  ����t$�@<��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh8�h�   h� ���V�  ����t���   ��t�MQ����^]� 3�^]� �U��Vh8�h�   h� ����  ����t���   ��t�MQ����^]� 3�^]� �U��Vh8�h�   h� �����  ����t'���   ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �U��Vh8�h�   h� ����  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h�   h� ���6�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h�   h� �����  ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh8�h�   h� ����  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h�   h� ���F�  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh8�h�   h� �����  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h�   h� ����  ����t,���   ��t"�E�M�U���$Q�MR�UQR����^]� 3�^]� ������������U��Vh8�h�   h� ���F�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h�   h� �����  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh8�h�   h� ����  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h�   h� ���V�  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h�   h� ����  ����tG���   ��t=�E(�MP���ĉ�M�H�M�H�M�H�M �H�M$�H�E�MPQ����^]�$ 3�^]�$ �U��Vh8�h�   h� ����  ����tN���   ��tD�E0�E(�MP�� ���\$��M�H�M�H�M�H�M �H�M$�H�E�MPQ����^]�, 3�^]�, ����������U��Vh8�h�   h� ����  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h   h� �����  ����t��   ��t�M�UQR����^]� 3�^]� �������������U��Vh8�h  h� ���v�  ����t#��  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh8�h  h� ���&�  ����t��  ��t�M�UQR����^]� 3�^]� �������������U��Vh8�h  h� �����  ����t��  ��t�M�UQR����^]� 3�^]� �������������U��Vh8�h  h� ����  ����t'��  ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �U��Vh8�h  h� ���6�  ����t#��  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh8�h  h� �����  ����t'��  ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �U��Vh8�h  h� ����  ����t��  ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h   h� ���F�  ����t��   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h$  h� �����  ����t#��$  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh8�h(  h� ����  ����t#��(  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh8�h,  h� ���V�  ����t3��,  ��t)�M$�U Q�MR�UQ�MR�UQ�MR�UQR����^]�  3�^]�  �����U��Vh8�h0  h� �����  ����t��0  ��t�MQ����^]� ��������U��Vh8�h4  h� ����  ����t��4  ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h8  h� ���f�  ����t��8  ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh8�h<  h� ����  ����t#��<  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh8�h@  h� �����  ����t#��@  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh8�hD  h� ���v�  ����t��D  ��t�M�UQ�MRQ����^]� U��Vh8�hH  h� ���6�  ����t��H  ��t�M�UQ�MRQ����^]� U���V��FT��u
���^��]� �V$�MjRP�E�M�P�M��E�����  ��t�+FT^����]� �����U���V��FX��u
���^��]� �V(�MjRP�E�M�P�M��E����F�  ��t�+FX^����]� �����U���V��F\��u
���^��]� �V,�MjRP�E�M�P�M��E������  ��t�+F\^����]� �����U���V��FL��u
���^��]� �V4�MjRP�E�M�P�M��E�Ĕ�E�������  ��t�+FL^����]� ��������������U���V��F<��u
���^��]� �V$�MjRP�E�M�P�M��E�̔�F�  ��t�+F<^����]� �����U���V��F@��u
���^��]� �V(�MjRP�E�M�P�M��E�̔���  ��t�+F@^����]� �����U���V��FD��u
���^��]� �V,�MjRP�E�M�P�M��E�̔��  ��t�+FD^����]� �����U���V��FP��u
���^��]� �V �MjRP�E�M�P�M��E����V�  ��t�+FP^����]� �����U���V��FH��u
���^��]� �V0�MjRP�E�M�P�M��E�Ĕ�E��������  ��t�+FH^����]� ��������������U���V��F8��u
���^��]� �V �MjRP�E�M�P�M��E�̔��  ��t�+F8^����]� �����U��E�@�M+A]� �������������U��E� �M+]� ���������������U��V�u���t�$��QP��Ѓ��    ^]���������̡$��H��@  hﾭ���Y����������U��E��t�$��QP��@  �Ѓ�]����������������U��$��H���  ]��������������U��$��H��  ]�������������̡$��H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW�Q0 ������u_^]Ã} tWj V��0 ��_������F�<�   ^]���U��$��ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW��/ ������u_^]�Wj V�0 ��_������F�<�   ^]�������������U��$��ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW�U/ ������u_^]�Wj V�0 ��_������F�<�   ^]�������������U��$��ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW��. ������u_^]�Wj V�/ ��_������F�<�   ^]�������������U��$��ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW�U. ������u_^]�Wj V�/ ��_������F�<�   ^]�������������U��M��t-�=<� t�y���A�uP�8/ ��]á$��P�Q�Ѓ�]��������U��M��t-�=<� t�y���A�uP��. ��]á$��P�Q�Ѓ�]��������U��$��H�U�R�Ѓ�]���������U��$��H�U�R�Ѓ�]���������U��$��ɋEt#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�- ������u_^]�Wj V��- ��_������F�<�   ^]���������U��$��ɋEtL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËMQ������]�������U��E��w�   �$���t�U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�", ������u_^]�Wj V��, ��_������F�<�   ^]����������U��E��w�   �$���t,�} �U�IR�URPt���   �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW�+ ������u_^]�Wj V�@, ��_������F�<�   ^]�������U��$��H�U�R�Ѓ�]���������U��$��H�U�R�Ѓ�]���������U��$��H�U�R�Ѓ�]���������U��$��H�U�R�Ѓ�]���������U��$��Hp�]��$��Hp�h   �҃�������������U��V�u���t�$��QpP�B�Ѓ��    ^]���������U��$��Pp�EP�EPQ�J�у�]� U��$��Pp�EP�EPQ�J�у�]� U��$��Pp�EP�EPQ�J�у�]� U��$��Pp�EPQ�J�у�]� ���̸   � ��������� ������������̃��� ����������� �������������U��$��H�QV�uV�҃���^]� ̸   � ��������3�� ����������̸   @� ��������3��  ����������̸   � ��������U��W�}��u3�_]� ��U�@@VR�Ћ���u^_]� �$��Q0�F�M���   PQW�ҋF��^_]� U��$��H0�U�AR�Ѓ���t
��ȋj��]� �������3�� ��������������������������̸   � ��������3�� �����������3�� �����������U��E� ����]� �������������̸   � ��������U��E� ����]� ��������������3�� �����������U��$��H���  ]��������������U��$��H���  ]��������������U��$��P�EP�EP�EP�EPQ���   �у�]� �����U��$��E�P�EP�E���\$�E�$PQ���   �у�]� �������������U��$��P�EP�EP�EPQ���   �у�]� ��������̡$��P���   Q�Ѓ�������������U��$��P�EP�EP�EPQ���   �у�]� ���������U��$��P�EP�EPQ���   �у�]� �������������U��$��H�U�ApR�Ѓ�]� �����U��$��P�EP�EPQ���  �у�]� �������������U��$��P�EP�EPQ���  �у�]� �������������U��$��P�EP�EPQ���  �у�]� �������������U��$��P�EP�EPQ���  �у�]� �������������U����   V�u��u3�^��]�Wh�   ��0���j P�t& ��R���E�P���ҡ$��P�B<�M��Ѕ��}t0j �M�QW�a�������u�$��B�P�M�Q�҃�_3�^��]ËE�M�Uh�   ��p�����0���P��t����MQWj	��P�����0���ǅ4����] �E��P�E�� �E�P� �E��P�E��P�E�� �E��Pǅx���p� ǅ|���pP�E��P�E��P�E��� �E� � �E�`� �E�П �E��� �E�0� �E�@� �E� � �EĀ� ��  �$����B�P�M�Q�҃�_��^��]����������U���   SV�u(3ۅ��]�u�$��H�A�UR�Ѓ�^3�[��]Ë$��Q�B<W�M3��Ѕ��'  ��  ���E�tq�MQ�M��il  WhД�M��{r��P�M��Rl  �u�Wj��U�R�E�P��\���Q�_?��  ��P��x���R�p  ��P�E�P��o  ��P�����  ���E�t�E� �� t�M�����pl  ��t��x�������]l  ��t��\�������Jl  ��t�M̃���:l  ��t�$��Q�J�E�P����у���t�M��l  �}� t"�U(�E$�M�R�UP�EQ�MRPQ���������U�R��  ����E$�M�UVP�Ej QRP����������$��Q�J�EP�у���_^[��]����������������U��E�M�UP�EQ�Mj RPQ������]�������������̋�`<����������̋�`L����������̋�`P����������̋�`����������̋�`����������̋�`$����������̋�`D����������̋�`T����������̋�`����������̋�`(����������̋�`H����������̋�`����������̋�`���������������P�P��P(�P �P�P@�P8�P0�PX�PP�PH����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX��������U��M�A8��   �IXV�AP�I@���I�AP�I(�AX�I ���I0���A@�I �A8�I(���IH����������Dz�u�؋��5�����^��]���W���A�IX�AP�I�A8�I�A�I@�AP�I@�U��A8�IX�]������IH�����I0�����e��	����ݝx����A�I(�U��A�I �U��AX�I �]��AP�I(�����IH�E����	���������I�������]��A8�I(�A@�I �����	�������I���E��e��I0�������]��E��e����]����e��ˋE��x������]������]��AH�I@�A0�IX�����]��AX�I�AH�I(�����]��A0�I(�A@�I�����]��AP�I0�AH�I8�����]��AH�I �AP�I�����]��A8�I�A0�I �   �����]��_^��]�������U��y0 ts��U�����Au���A�Z����Au�B�Y�A�Z����Au�B�Y�A�����z��Y�A �Z����z�B�Y �A(�Z����zZ�B�Y(]� �E��Q�P�Q�P�Q �P�Q$�P�Q(�@�A,�Q�A��Q �A�A$�Q�Q(�A�A,�Q�A�A0   ]� U��y0 tL��E�A�A �A�A(�A�������������X�X�A� �A �`�A(�`�E����X�X]� ��E����������P���P�E����X�X]� ��̋�3ɉ�H�H�H�V��V�����FP����3����F�F^��3���A�A�A����A�`�
�@�b�	���B�a�������U����   ��UV���q�U�W3��<��M��}���  ��S�]�k  ��؋�U��M�U��U�@�����@�U��@�B�@�������@���@�G�>��w����U���  �w������݃��B��   �U������ɋP��R�э����]��B���B�P���R���U����E������]��E��M��E������������]��E����E����E��E��]����E��]����E��]��]����U��E��U�����B���B���U������������]��E����E����������E������E��E��]����E��]����E��]����U��E��]���R�э�������B���B�P���R���U����E��������]��E����E����������E������E��E��]��E��]����E��]��U��E��]�����B���B���U����E��������]��E����E����������E������E��E��]��E��]����E��]��E��U��`�����E�U���������;���   �ލ�+���͋�@����������]��@���]��@���U������M������]��E��E����E��������]��E������������E��E��]��E��E��]����E��]��E��U�u�������������������������������M���Q�ʍU��R���[�[�kh����E�KH��P�E��SL��H�щKP�P�ST�H�KX�P�������S\z^�E�����������zP���CP�����CX���CH���CX�������cH���[�[ �[(�C(�KP�C �KX���C�KX�C(�KH���CH�K �\���E���������za�CX�����CP�����cH�CH���CP�������[���[ �[(�CP�K(�C �KX���C�KX�CH�K(���C �KH�C�KP�����[0�[8�[@�[�CP�����CX�����KH�CX�����cP���[0�[8�[@�C8�KX�C@�KP���C@�KH�CX�K0���CP�K0�C8�KH�����[�[ �[(��$���SP������E��U�   �����}��M�����م�~�A8����u��1���U�@���K�I��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�@�K@���CX�H�D��@�����U���]��C���@�K0���CH�H���C ��C�@�K8���@�KP���C(��C�C@�H���CX�H3������U��x  �A������܃��E����E   �E�
���������ɋE������׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H�E������������������������������E����]��E��]����]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H�E��������]������M������������������������]��E��]��E��]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H���]������M������������������������]��E�Eȃ��]���E����]ȃE׃m����@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H���]������M������������������������U��E��]��E��U�������E������������;���   �P�U��+ЉU�
���������ʋE���׋��U�@���K��@�K0���CH�H���]�� �K �C�@�K8���@�KP���]�� �K(�C�C@�H���CX�H�   E)E���]����E��������������������M����������]��E��E��U�����[������_��^��]� ��[��_��^���؋�]� �����������h@�Ph_� ��  ���������������h@�jh_� �϶  ����uË@����U��V�u�> t/h@�jh_� 裶  ����t��U�M�@R�Ѓ��    ^]���U��Vh@�jh_� ���i�  ����t�@��t�MQ����^]� 3�^]� �������U��Vh@�jh_� ���)�  ����t�@��t�MQ����^]� 3�^]� �������U��Vh@�jh_� ����  ����t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh@�jh_� ��虵  ����t�@��t�MQ����^]� 3�^]� �������U��Vh@�j h_� ���Y�  ����t�@ ��t�MQ����^]� 3�^]� �������U��Vh@�j$h_� ����  ����t�@$��t�MQ����^]� 2�^]� �������Vh@�j(h_� ���ܴ  ����t�@(��t��^��3�^������Vh@�j,h_� ��謴  ����t�@,��t��^��3�^������U��Vh@�j0h_� ���y�  ����t�@0��t�MQ����^]� 3�^]� �������U��Vh@�j4h_� ���9�  ����t�@4��t�M�UQR����^]� ���^]� ��Vh@�j8h_� �����  ����t�@8��t��^��3�^������U��Vh@�j<h_� ���ɳ  ����t�@<��t�MQ����^]� ��������������U��Vh@�j@h_� ��艳  ����t�@@��t�MQ����^]� ��������������U��Vh@�jDh_� ���I�  ����t�@D��t�MQ����^]� 3�^]� �������U��Vh@�jHh_� ���	�  ����t�@H��t�MQ����^]� ��������������Vh@�jLh_� ���̲  ����t�@L��t��^��3�^������Vh@�jPh_� ��蜲  ����t�@P��t��^��3�^������Vh@�jTh_� ���l�  ����t�@T��t��^��^��������Vh@�jXh_� ���<�  ����t�@X��t��^��^��������Vh@�j\h_� ����  ����t�@\��t��^��^��������U��Vh@�j`h_� ���ٱ  ����t�@`��t�M�UQR����^]� 3�^]� ���U��Vh@�jdh_� ��虱  ����t�@d��t�M�UQR����^]� 3�^]� ���U��Vh@�jhh_� ���Y�  ����t�@h��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh@�jlh_� ���	�  ����t�@l��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh@�jph_� ��蹰  ����t�@p��t�M�UQR����^]� 3�^]� ���U��Vh@�jth_� ���y�  ����t�@t��t�M�UQR����^]� 3�^]� ���U��Vh@�jxh_� ���9�  ����t�@x��t�M�UQR����^]� 3�^]� ���U��Vh@�j|h_� �����  ����t�@|��t�MQ����^]� 3�^]� �������U��Vh@�h�   h_� ��趯  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh@�h�   h_� ���f�  ����t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh@�h�   h_� ����  ����t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh@�h�   h_� ��覮  ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U���|��A�����U����U����U��  S�V�E��EW�����������   ���������U�r�z�
�R;��4v���4��I�$ȍ��F�R�a���F�a�uB�!�]��B�a�U��B�a�U������������]��E����E����������E��������E��G��$ȍ��]��B�a�U��B�a�U������������]��E����E����������E��������E��������m�������_�U�^��[�U����U�������������������� ����������D�Ez���P�P���]� �������E�����E����X�M��X��]� �������U���@�H��A�������E�    ���]����]��]��ؔ�������]����]��]���   �	S�]VW�M��E����������t[��%�����E�M�����@��P������F�@��R�M������~���Q�M������v;�t�v��P�M������M����m��M�u�_^[�M�UQR�M��A�����]� ����������̋Q3���|�	��t��~�    t������u��3�������U��QV�u;��}�	���    u����;�|���^]� +ƃ�^]� �������U��VW�}��|-�1��t'�Q3���~�΍I �1�������;�t����;�|���_^]� �������������̋Q3���~%V�1�d$ ���   @u�����t������u�^�̋QV3���~�	�d$ ����Шt������u��^�������U��Q3�9A~��I ��$��������;A|�Q��~[SVW�   3ۋ���x5��%���;��E���}$��������%���;E�u�
   ���;q|݋Q���G���;�|�_^[��]�������U��	����%�����E��   @t����������wg�$��� �E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� T� j� }� �� �� ����U����S��V������   @Wt���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V��V�g����FP�^���3����F�F^��U��SV��WV�B����^S�9����E3���;ǉ~�~t_�$��Q���   h����jIP�у�;ǉt9�}��t;�$��B���   h����    jNQ�҃����uV�������_^3�[]� �E�~_�F^�   []� ����������U��SV��WV�����^S�����}3Ƀ�;��N�N��   9��   �G;���   �$��Q���  h����jlP�у����t=� t@�G��t9�$��Jh����    ���  jqR�Ѓ����u���]���_^3�[]� �O�N�G�Q��    R�F�QP�L  �����t�N�WP��QPR�xL  ��_^�   []� ���������U��SV��WV�����~W����3Ƀ�9M�N�N��   �E;���   ��    �$��H���  h��h�   S�҃����t=�} tH�E��tA�$��Q���  h����h�   P�у����u���b���_^3�[]� �U�V�,�F   �$��H���  h��h�   j�҃����t��E�M�F�PSPQ�qK  �E����t!�V�?�W�RWP�UK  ��_^�   []� ��M�_^�   []� ���U��Q2���~CS�]V�1W������������;�u��   @u�����u3���   ��
���u�_^[��]� �����������U��S�]V��3�W�~���F�F�C;CV��   �����W�����3��F�F�$��Q���   h��jIj�Ѓ������   �$��Q���   h��jNj�Ѓ����uV������_��^[]� ��F   �F   ����K�H�C��B�_��^�   []� �@���W�:���3��F�F�$��B���   h��jIj�у����t[�$��B���   h��jNj�у�����\�����F   �F   ����S�Q��K�H��C�B��   _��^[]� �����������U��3�V���F�F�F�EP�������^]� �������������U��EVP���������^]� ���������̡$��HL���   ��U��$��H@�AV�u�R�Ѓ��    ^]�������������̡$��HL�������U��$��H@�AV�u�R�Ѓ��    ^]�������������̡$��PL���   Q�Ѓ�������������U��$��PL�EP�EPQ���   �у�]� �������������U��$�V��HL���   V�҃���u�$��U�HL���   j RV�Ѓ�^]� �$����   �ȋBP�Ћ$����   �MP�BH��^]� �����̡$��PL��(  Q�Ѓ�������������U��$��PL�EP�EPQ��,  �у�]� ������������̡$��HL�Q�����U��$��H@�AV�u�R�Ѓ��    ^]��������������U��$��PL�E�R��VPQ�M�Q�ҋu��P���ň  �M��݈  ��^��]� ����U��$��PL�EPQ���   �у�]� �U��$��PL�EP�EPQ�J�у�]� �$��PL�BQ�Ѓ���������������̡$��PL�BQ�Ѓ���������������̡$��PL�BQ�Ѓ����������������U��$��PL�EP�EP�EPQ�J �у�]� ������������U��$��PL�EPQ��4  �у�]� �U��$��PL�EP�EP�EPQ�J$�у�]� ������������U��$��PL�EP�EP�EP�EPQ�J(�у�]� �������̡$��PL�B,Q�Ѓ���������������̡$��PL�B0Q�Ѓ����������������U��$��PL�EP�EPQ��  �у�]� ������������̡$��PL���   Q�Ѓ�������������U��$��PL�E��  ��VPQ�M�Q�ҋu��P��袆  �M�躆  ��^��]� ̡$��PL�B4Q�Ѓ���������������̡$��PL�B8j Q�Ѓ��������������U��$��PL���   ]��������������U��$��PL���   ]��������������U��$��PL���   ]��������������U��$��PL���   ]��������������U��$��PL���   ]��������������U��$��PL���   ]��������������U��$��PL���   ]��������������U��$��PL���   ]��������������U��$��PL���   ]��������������U��$��PL�EPQ�J<�у�]� ���̡$��PL�BQ��Y�U��$��PL�EP�EPQ�J@�у�]� U��$��PL�Ej PQ�JD�у�]� ��U��$��PL�Ej PQ�JH�у�]� ��U��$��PL�EjPQ�JD�у�]� ��U��$��PL�EjPQ�JH�у�]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}�蔘  W�M�Q�U�R���4�  ���M������  ��t�$����   ��U�R�Ѓ�_^3�[��]Ë$����   �J8�E�P�ы$������   ��M�Q�҃�_��^[��]��������������U���$3�V�E��E�E��P�M��E�   �E�   �E��  �ޗ  j�M�Q�U�R��蝺  �M��E�  �$����   ��U�R�Ѓ�^��]�����������U���$�$��UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��Z�  j�E�P�M�Q����  �M����  �$����   ��M�Q�҃�_^��]� ��U���$�$��UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��ږ  j�E�P�M�Q��虹  �M��A�  �$����   ��M�Q�҃�_^��]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��t�  W�M�Q�U�R����  ���M����׈  ��t+�u����@  �$����   ��U�R�Ѓ�_��^[��]� �$����   �JL�E�P�ыu��P���EA  �$����   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}�贕  W�M�Q�U�R���T�  ���M�����  ��t+�u���@  �$����   ��U�R�Ѓ�_��^[��]� �$����   �JL�E�P�ыu��P���@  �$����   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}����  W�M�Q�U�R��蔷  ���M����W�  _^��[t�$����   ��U�R�������]Ë$����   �J<�E�P���]��$����   ��M�Q���E�����]���������������U���$SVW3��E��P�M��}܉}��E��  �}��}��D�  W�M�Q�U�R����  ���M���视  ��t�$����   ��U�R�Ѓ�_^3�[��]Ë$����   �J8�E�P�ы$������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}�蔓  W�M�Q�U�R���4�  ���M������  ��t-��u�$�����   ���^�U�R�Ѓ�_��^[��]� �$����   �JP�E�P�ы�u�H��P�@�N�$��V���   �
�F�E�P�у�_��^[��]� �����̡$��PL���   Q��Y��������������U��$��PL�E���   ��jPQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U��$��PL�E���   ��j PQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���$SVW3��E��P�M��}܉}��E��  �}��}���  W�M�Q�U�R��褴  ���M����g�  ��t-��u�$�����   ���^�U�R�Ѓ�_��^[��]� �$����   �JP�E�P�ы�u�H��P�@�N�$��V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��4�  W�M�Q�U�R���Գ  ���M���藃  ��t-��u�$�����   ���^�U�R�Ѓ�_��^[��]� �$����   �JP�E�P�ы�u�H��P�@�N�$��V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��d�  W�M�Q�U�R����  ���M����ǂ  ��t-��u�$�����   ���^�U�R�Ѓ�_��^[��]� �$����   �JP�E�P�ы�u�H��P�@�N�$��V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}�蔏  W�M�Q�U�R���4�  ���M������  ��t�$����   ��U�R�Ѓ�_^3�[��]Ë$����   �J8�E�P�ы$������   ��M�Q�҃�_��^[��]��������������U����E3�V�]�E��E��E��P�M�E�   �E��  �ߎ  j�M�Q�UR��螱  �M�F�  �$����   ��U�R�Ѓ�^��]� ���������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��o�  j�U�R�E�P���.�  �M��ր  �$����   �
�E�P�у�^��]� ��������U���$�$��UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}���  j�E�P�M�Q��詰  �M��Q�  �$����   ��M�Q�҃�_^��]� ��U���$�$��UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��j�  j�E�P�M�Q���)�  �M���  �$����   ��M�Q�҃�_^��]� ��U���$�$��UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}���  j�E�P�M�Q��詯  �M��Q  �$����   ��M�Q�҃�_^��]� ��U���$�$��UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��j�  j�E�P�M�Q���)�  �M���~  �$����   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E����  j�U�R�E�P��辮  �M��f~  �$����   �
�E�P�у�^��]� ��������U���$SVW3��E��P�M��}܉}��E��  �}��}�蔋  W�M�Q�U�R���4�  ���M�����}  ��t-��u�$�����   ���^�U�R�Ѓ�_��^[��]� �$����   �JP�E�P�ы�u�H��P�@�N�$��V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��Ċ  W�M�Q�U�R���d�  ���M����'}  ��t�$����   ��U�R�Ѓ�_^3�[��]Ë$����   �J8�E�P�ы$������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}���  W�M�Q�U�R��贬  ���M����w|  ��t�$����   ��U�R�Ѓ�_^3�[��]Ë$����   �J8�E�P�ы$������   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ����U���$�$��UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��*�  j�E�P�M�Q����  �M��{  �$����   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E�迈  j�U�R�E�P���~�  �M��&{  �$����   �
�E�P�у�^��]� ��������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��O�  j�U�R�E�P����  �M��z  �$����   �
�E�P�у�^��]� ��������U��$��H���   ]��������������U��$��H���   ]�������������̡$��H���   ��$��H���   ��U��$��H���   V�u�R�Ѓ��    ^]�����������U��$��H���   ]��������������U��$��HL�QV�ҋ���u^]á$��H�U�ER�UP���  RV�Ѓ���u�$��Q@�BV�Ѓ�3���^]����������U��$��H�U�E���  R�U�� P�ERP�у�]������U��$��H���   ]��������������U��$��H�U �ER�UP�ER�UP�ER�UP���   R�Ѓ�]������������̡$��PL�BLQ�Ѓ���������������̡$��PL�BPQ�Ѓ����������������U��$��PL�EP�EPQ�JT�у�]� U��$��PL�EPQ��  �у�]� �U��$��PL�EPQ���   �у�]� ̡$��PL�BXQ�Ѓ����������������U��$��PL�EP�EP�EPQ�J\�у�]� ������������U���4�$�SV��HL�QW�ҋ�3�;��}��x  �M��p  �$��E�EԋE�]Љ]؉]܉]�]��}̋Q�R0Ph]  �M��ҡ$����   �BSSW���Ѕ���   �$��QL�BW�Ћ���;���   ��    �$����   �B(���ЍM�Qh�   ���u��zW  ������   �M�;���   �$����   ���   S��;�tm�$����   �ȋB<V�Ћ$����   ���   �E�P�у�;�t�$��B@�HV�у�;����\����}��M��Qk  �M���o  ��_^[��]� �}��$��B@�HW�ы$����   ���   �M�Q�҃��M��	k  �M��o  _^3�[��]� �����̡$��PL�B`Q�Ѓ���������������̡$��PL�BdQ�Ѓ����������������U��$��PL�EPQ�Jh�у�]� ���̡$��PL��D  Q�Ѓ������������̡$��PL�BlQ�Ѓ����������������U��$��PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U$�EV�Eh�� h�� h�� h�� R�Q�U R�UR�UR�U���A�$�5$��vLRP���   Q�Ѓ�4^]�  ������̡$��PL���   Q�Ѓ�������������U��$��PL�EP�EP�EPQ��   �у�]� ���������U��$��PL��H  ]�������������̡$��PL��L  ��U��$��PL��P  ]��������������U��$��PL��T  ]��������������U��$��PL�EP�EP�EP�EP�EPQ���   �у�]� �U��$��PL�EP�EP�EPQ���   �у�]� ���������U��$��PL�EP�EP�EP�EPQ��   �у�]� �����U��$��HL���   ]��������������U��$��HL���   ]��������������U��$��HL���   ]�������������̡$��HL��  ��$��HL��@  ��hT�Ph^� � �  ���������������U��VhT�j\h^� �����  ����t�@\��t
�MQV�Ѓ�^]� ������������U��� �$�V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ};��E�t`;�t\�$��QLjP���   ���ЋM��U�Rh=���M�}��cR  ���$����   ���   �U�R�Ѓ��M��u��f  ��_^��]Ë$����   ���   �E�P�у��M��u��nf  _�   ^��]����U��� �$�V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ};��E�t`;�t\�$��QLjP���   ���ЋM��U�Rh<���M�}��Q  ���$����   ���   �U�R�Ѓ��M��u���e  ��_^��]Ë$����   ���   �E�P�у��M��u��e  _�   ^��]����U��$��E�PH�B���$Q�Ѓ�]� ���������������U��$��PH�EPQ���   �у�]� �U��$��PH�EPQ���  �у�]� �U��$��PH�EPQ���  �у�]� �U��$��PH�EP�EPQ��  �у�]� �������������U��$��PH�EP�EPQ��  �у�]� ������������̡$��PH���  Q�Ѓ�������������U��$��PH�EPQ���  �у�]� ̡$��PH���   j Q�Ѓ�����������U��$��PH�EPj Q���   �у�]� ��������������̡$��PH���   jQ�Ѓ�����������U��$��PH�EPjQ���   �у�]� ��������������̡$��PH���   jQ�Ѓ����������U��$��PH�EPjQ���   �у�]� ���������������U��$��PH�EP�EPQ���   �у�]� �������������U��$��PH�EP�EPQ���   �у�]� ������������̡$��PH���   Q�Ѓ�������������U��$��PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP����  ������t�E�$��QH���   PVW�у���_^]� �����U��EVW���MPQ��  ������t�M�$��BH���   QVW�҃���_^]� ̡$��PH���   Q�Ѓ������������̡$��PH���   Q�Ѓ�������������U��$��PH�EPQ���   �у�]� �U��$��PH�EPQ���   �у�]� �U��$��PH�EP�EPQ��8  �у�]� �������������U��$��PH�EP�EPQ��   �у�]� ������������̡$��PH���  Q�Ѓ������������̡$��PH���  Q�Ѓ������������̡$��PH���  Q�Ѓ������������̡$��PH��  Q�Ѓ������������̡$��PH��  Q�Ѓ�������������U��$��PH�EP�EPQ��  �у�]� �������������U��$��PH�EP�EP�EPQ��   �у�]� ���������U��$��PH�EP�EP�EP�EPQ��|  �у�]� �����U��$��PH�EPQ��  �у�]� ̡$��PH��T  Q�Ѓ�������������U��$��PH�EP�EPQ��  �у�]� �������������U��$��PH�EPQ��8  �у�]� �U��$��PH�EPQ��<  �у�]� �U��$��PH�EPQ��@  �у�]� �U��$��PH�EP�EP�EPQ��D  �у�]� ��������̡$��PH��L  Q��Y��������������U��$��PH�EPQ��H  �у�]� ̡$�V��H@�Q,WV�ҋ$��Q��j �ȋ��   h�  �Ћ$��QH�����   h�  V�Ѓ���
��t_3�^Ë�_^�̡$��P@�B,Q�Ћ$��Q��j �ȋ��   h�  �������U��$��E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U��$��E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U��$��PH�EP�EP�EPQ��   �у�]� ��������̡$��HH��  ��U��$��HH��  ]��������������U��$��E�PH��$  ���$Q�Ѓ�]� �����������̡$��PH��(  Q�Ѓ�������������U��$��PH�EP�EPQ��,  �у�]� �������������U��$��E�PH�EP�E���$PQ��0  �у�]� ���̡$��PH���  Q�Ѓ������������̡$��PH��4  Q�Ѓ������������̋��     �������̡$��PH���|  jP�у���������U��$��UV��HH��x  R��3Ƀ������^��]� ��̡$��PH���|  j P�у��������̡$��PH��P  Q�Ѓ������������̡$��PH��T  Q�Ѓ������������̡$��PH��X  Q�Ѓ�������������U��$��PH��Q��\  �E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����̡$��PH��`  Q�Ѓ�������������U��$��PH�EPQ��d  �у�]� �U��$��E�PH��h  ���$Q�Ѓ�]� ������������U��$��E�PH��t  ���$Q�Ѓ�]� ������������U��$��E�PH��l  ���$Q�Ѓ�]� ������������U��$��PH�EPQ��p  �у�]� �U��$��PH�EP�EP�EP�EPQ���  �у�]� �����U��$��PH�EP�EP�EP�EP�EP�EPQ���  �у�]� �������������U��$��E�HH�U �ER�UP�E���$R�UP���   R�Ѓ�]������������U��U�E�$��HH�E���   R�U���$P�ERP�у�]����������������U���E�M������  �M;�|�M;�~��]�����������U��$��PH�E���   Q�MPQ�҃�]� ������������̡$��PH���   Q��Y�������������̡$��PH���   Q�Ѓ������������̡$��PH���   Q��Y��������������U��$��PH�EP�EPQ���   �у�]� �������������U��$��PH�EP�EP�EP�EP�EPQ���  �у�]� ̡$��PH��t  Q��Y�������������̋��  ��@    �� ��$��Pl�A�JP��Y��������U��$�V��Hl�V�AR�ЋE����u
�   ^]� �$��Ql�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uË$��QlP�B�Ѓ�������U��$��Pl�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U��U�E�$��HH�ER�U���$P���  R�Ѓ�]����U��$��HH���  ]��������������U��$��HH���  ]��������������U��U0�E(�$��HH�E$R�U ���$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�,]������������U��$��HH���  ]��������������U��$��E�PH�EP���$Q���  �у�]� ��������U���SV���V  �؅ۉ]���   �} ��   �$��HH��p  j h�  V�҃����E�u
^��[��]� �MW3��}��V  ����   �]��I �E�P�M�Q�MW�OW  ��tc�u�;u�[�I ������u�E�������L�;Ht-�$��Bl�S�@����QR�ЋD������t	�M�P�3V  ��;u�~��}��M���}���U  ;��r����]�_^��[��]� ^3�[��]� ����������U����$�SV�ًHH��p  j h�  S�]��ҋ�����u
^3�[��]� �E��u�$��HH���  �'��u�$��HH���  ���uš$��HH���  S�ҋȃ��ɉEt�W��U  �$��HH���   h�  S3��҃����  ���_�u����    �$��Hl�U�B�IWP�ы�������   �$��F�J\�UP�A,R�Ѓ���t�K�Q�M��T  �$��F�J\�UP�A,R�Ѓ���t�K�Q�M�T  �E��;Pt&�F�$��Q\�J,P�EP�у���t	�MS�T  �$��v�B\�M�P,VQ�҃���t�M�CP�cT  �$��QH�E����   �E�h�  P�����у�;�����_^�   [��]� ������U��$��HH���   ]�������������̡$��PH���   Q��Y��������������U��$��HH���  ]��������������U��$���P���   V�uW�}���$V�����E������At���E������z����؋$��Q�B,���$V����_^]����������������U���0��$��U�V�u�U��]�W�P�}���   �E�PV�M�Q����� �@�@�E�����E��Au�����������z���������������z�����������Au������������z)���١$��]��ɋ��]��]��P�RH�E�PV��_^��]���������Au������������������U��$��HH�]��U��$��H@�AV�u�R�Ѓ��    ^]�������������̡$��HH�h�  �҃�������������U��$��H@�AV�u�R�Ѓ��    ^]��������������U��$��HH�Vh  �ҋ�������   �EPh�  ��  ����t]�$��QHj P���   V�ЋMQh(  �Ƶ  ����t3�$��JH���   j PV�ҡ$����   �B��j j���Ћ�^]á$��H@�QV�҃�3�^]�������U��$��H@�AV�u�R�Ѓ��    ^]��������������U��$��HH�Vh�  �ҋ�����u^]á$��HH�U�E��  RPV�у���u�$��B@�HV�у�3���^]�������U��$��H@�AV�u�R�Ѓ��    ^]��������������U��$��HH�I]�����������������U��$��H@�AV�u�R�Ѓ��    ^]��������������U��$��PH�EPQ���  �у�]� �U��$��PH�EPQ���  �у�]� ̡$��PH���  Q�Ѓ�������������U��$��HH���  ]��������������U��$��E�HH�U0�E,R�U(P�E$R�U P�ER�U���\$�E�$P��P  R�Ѓ�,]������������̡$��PH���  Q�Ѓ�������������U��$��PH�EP�EPQ���  �у�]� ������������̡$��PH��  Q�Ѓ�������������U��$��PH�EP�EP�EPQ���  �у�]� ��������̡$��PH���  Q�Ѓ������������̡$��PH���  Q�Ѓ�������������U��$��PH�EPQ��  �у�]� �U��$��PH�EPQ��  �у�]� ̋������������������������������̡$��HH���  ��U��$��HH���  ]��������������U��$��PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ���������U��$��PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ��������̡$��PH��,  Q�Ѓ�������������U��$��PH�EPQ��X  �у�]� ̡$��PH��\  Q�Ѓ�������������U��$��HH��0  ]��������������U��$���W���HH���   j h�  W�҃��} u�   _��]� Vh�  �o�  ��������   �$��HH���   j VW�҃��M��O  �$��P�E�R0Ph�  �M����E�$��P�B,���$h�  �M��Ћ$��Q@�J(j �E�PV�у��M��O  ^�   _��]� ^3�_��]� �����U��S�]�; VW��u7�$��U�HH���   RW�Ѓ���u�$��QH���   jW�Ѓ���t�   �����   �$��QH���   W�Ѓ��} u(�$��E�QH�M���  P�ESQ�MPQW�҃��B�u��t;�$��U�HH�ER�USP���  VRW�Ћ$����   �B(�����Ћ���uŃ; u�$��QH���   W�Ѓ���t3���   ���Wu1�$��QH���   �Ћ$��E�QH���   PW�у�_^[]� �$��BH���   �у��} u0�$��M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� �$��QH�h  �Ћ؃���u_^[]� �$����   �u�Bx���Ћ$����   P�B|���Ѕ�tU�$��E�QH�MP�Ej Q���  VPW�у���t�$����   �ȋBHS�Ћ$����   �B(���Ћ���u�_^��[]� ��������������U��E��V��u�$��HH���  �'��u�$��HH���  ���u�$��HH���  V�҃���u3�^]� P�EP���>���^]� ���������U���D�$��HH���   S�]VWh�  S�ҋ�$��HH���   3�Wh�  S�u܉}��҃�;��E�}�}��}��p
  �$����   �B����=�  �$��  �QH���   Wh:  S�Ћ$��QH�E����   h�  S�Ћ$��QHW�����   h�  S�uԉ}��Ћ$��QH�E苂  S�Ћ$��QH�EЋ��  S�Ѓ�(���E��E�,��}   �M���M�MЅ�tMj�W�P������t@�@�Ẽ|� �4�~����%�������;�u/���o���;E�~�E؋��0���E���E�;Pu�E���E��E���;}�|��}� tv�u�j S���h�  ����  ���Y�  ��tV�����  �}�;�uK�$��H���  �4�h0���h�  V�҃����E��k  �M�PVP�
�  P��  ����}ܡ$��H���  �4�h0���h�  V�҃����E��   �M�3�;�t;�tVQP��  ���E�;�~-�$��Qh0���h�  P���   �Ѓ�;ǉE���  �$��E��QH��  j�PS�у�����  �u�;�tjS���J�  ����  ���[�  �E���}�$��BH���   Wh�  S�у�3�9}ԉE�}���  �}���}ȋMЅ��p  �U�j�R�X�������\  �M̍@�|� ���]�~����%�������9E��  ���;����E�3�3�9C�E܉M���   ��I �����������t{�]��}������������ϋ9�<��}����҉��y�]��|��]������z�<��y�]��|��]������z�<��I�}��]������M��}ȃ��������M؃�;K�M��b������E��O  �+U�j��PR�M��f  �M�v���E�3�+��U��E����	��$    ���E�;E���   �}� �U����E�t6�U�@�U�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�M��E�;]؍@�E��Ћ��P�Q�P�Q�P�Q�P�Q�@�A}c�UȋE�9�uX�ȋL�����������w4�$�x	�U����4�"�M����t��U����t�
�M����t�M���;]�|��E�����;]؉M������U�;U��  �U�R�ь���E�P�Ȍ���M�Q迌����_^3�[��]Ë�M�3�;G�Å���   �E�v�ЋW��R�ы��Q�P�Q�P�Q�P�Q�P�I�H�O��I�M�ы�P�Q�P�Q���ۉP�Q�P�Q�P�I�H��@�E�ЋU�Lv�ʋ��P�Q�P�Q�P�Q�P�Q�@�At8�G�U�@�ʋU�Lv	�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��w��U��@�ʋU���v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��w��U����@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�7����t?�G�U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�w�����O�E�����;EԉE��}�������U�R觊���E�P螊�����$  ���   �B����=  �  �$��QH���   j h(  S�Ћ$��QH�����   h(  S�ЋЃ�3��҉U�~#���ǅ�t�|� t�4N��tN���;�|�u��u܋$��Q���  �4v�h0���hK  V�Ѓ����E���   �M��t��tVQP��  ���u؋$��Q���  �h0���hP  V�Ѓ����E�tP��t��tVWP���  ���M����+$��RH��PQ�E���   S�Ѓ���u�M�Q�\����U�R�S�����_^3�[��]á$��HH���   j h�  S�҉E��$��HH���   j h(  S��3�3���3�9]؉E��}ĉ]��N  �U���    �څ��+  ���E�    ��   �U�<��v��   ����U��:��\:�Y�\:�Y�\:׉Y�Z�Y�R�Q�U��\�E��Y�\�T���Y�Z�Y�Z�Y�Z�Y�R�]��Q�U�����������;�|��}ă|� �w   �U��Eԍ8�I�ʋU�v���A�B�A�B�A�B�A�B�I�J�E���ЋE���v�Ћ��A�B�A�B�A�B�A�B�I�J�U���<ډ}ă�;]؉]�������M�3�3�;�~"�U����$    �d$ �t���   ��;�|�U�R�u������E�P�i�����_^�   [��]Ë�������������U��U��t�M��t�E��tPRQ�P�  ��]������������U��V��V� ��$��Hl�AR�Ѓ��Et	V�$�������^]� ����������U��$��P�EP�EP�EPQ�J�у�]� �����������̡$�V��H�QV�ҡ$��H$�QDV�҃���^�����������U��$�V��H�QV�ҡ$��H$�QDV�ҡ$��U�H$�AdRV�Ѓ���^]� ��U��$�V��H�QV�ҡ$��H$�QDV�ҡ$��U�H$�ARV�Ѓ���^]� ��U��$�V��H�QV�ҡ$��H$�QDV�ҡ$��H$�U�ALVR�Ѓ���^]� �̡$�V��H$�QHV�ҡ$��H�QV�҃�^�������������U��$��P$�EPQ�JL�у�]� ����U��$��P$�R]�����������������U��$��P$�Rl]����������������̡$��P$�Bp����̡$��P$�BQ�Ѓ����������������U��$��P$��VWQ�J�E�P�ы$��u���B�HV�ы$��B�HVW�ы$��B�P�M�Q�҃�_��^��]� ���U��$��P$�EPQ�J�у�]� ����U��$��P$��VWQ�J �E�P�ы$��u���B�HV�ы$��B$�HDV�ы$��B$�HLVW�ы$��B$�PH�M�Q�ҡ$��H�A�U�R�Ѓ� _��^��]� ���U��$��P$��VWQ�J$�E�P�ы$��u���B�HV�ы$��B$�HDV�ы$��B$�HLVW�ы$��B$�PH�M�Q�ҡ$��H�A�U�R�Ѓ� _��^��]� ���U���V�uV�E�P�l������e����$��Q$�JH�E�P�ы$��B�P�M�Q�҃���^��]� ����̡$��P$�B(Q��Yá$��P$�BhQ��Y�U��$��P$�EPQ�J,�у�]� ����U��$��P$�EPQ�J0�у�]� ����U��$��P$�EPQ�J4�у�]� ����U��$��P$�EPQ�J8�у�]� ����U��$��UV��H$�ALVR�Ѓ���^]� ��������������U��$��H�QV�uV�ҡ$��H$�QDV�ҡ$��H$�U�ALVR�Ћ$��E�Q$�J@PV�у���^]�U��$��UV��H$�A@RV�Ѓ���^]� ��������������U��$��P$�EPQ�J<�у�]� ����U��$��P$�EPQ�J<�у������]� �������������U��$��P$�EP�EPQ�JP�у�]� U��$��P$�EPQ�JT�у�]� ���̡$��H$�QX�����U��$��H$�A\]�����������������U��$��P$�EP�EP�EPQ�J`�у�]� �����������̡$��H(�������U��$��H(�AV�u�R�Ѓ��    ^]��������������U��$��P(�R]����������������̡$��P(�B�����U��$��P(�R]�����������������U��$��P(�R]�����������������U��$��P(�R ]�����������������U��$��P(�E�RjP�EP��]� ��U��$��P(�E�R$P�EP�EP��]� �$��P(�B(����̡$��P(�B,����̡$��P(�B0�����U��$��P(�R4]�����������������U��$��P(�RX]�����������������U��$��P(�R\]�����������������U��$��P(�R`]�����������������U��$��P(�Rd]�����������������U��$��P(�Rh]�����������������U��$��P(�Rx]�����������������U��$��P(�Rl]�����������������U��$��P(�Rt]�����������������U��$��P(�Rp]�����������������U��$��P(�BpVW�}W���Ѕ�t:�$��Q(�Rp�GP���҅�t"�$��P(�Bp��W���Ѕ�t_�   ^]� _3�^]� ��U��$��P(�BtVW�}W���Ѕ�t:�$��Q(�Rt�GP���҅�t"�$��P(�Bt��W���Ѕ�t_�   ^]� _3�^]� ��U��VW�}W���0�����t8�GP���!�����t)�OQ��������t��$W��������t_�   ^]� _3�^]� ������������U��VW�}W���0�����t8�GP���!�����t)�O0Q��������t��HW��������t_�   ^]� _3�^]� ������������U����$��E�    �E�    �P(�RhV�E�P���҅���   �E���uG�$��H�A�U�R�Ћ$��Q�E�RP�M�Q�ҡ$��H�A�U�R�Ѓ��   ^��]� �$��Qhh�h`  P���   �Ћ$������E��Q(u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P�|����3�^��]� �M��U�j ���Q�MR�����E�P��{�����   ^��]� �������������U��$���V��H�A�U�R�Ѓ��M�Q��������^u�$��B�P�M�Q�҃�3���]� �$��H$�E�I�U�RP�ы$��B�P�M�Q�҃��   ��]� �U��Q�$��P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U��$��P(�R8]�����������������U��$��P(�R<]�����������������U��$��P(�R@]�����������������U��$��P(�RD]�����������������U��$��P(�RH]�����������������U��$��P(�E�R|P�EP��]� ����U��$��P(�RL]�����������������U��$��E�P(�BT���$��]� ���U��$��E�P(�BPQ�$��]� ����̡$��H(�Q�����U��$��H(�AV�u�R�Ѓ��    ^]��������������U��$��P(���   ]��������������U��$��H(�A]����������������̡$��H,�Q,����̡$��P,�B4�����U��$��H,�A0V�u�R�Ѓ��    ^]�������������̡$��P,�B8�����U��$��P,�R<��VW�E�P�ҋu���$��H�QV�ҡ$��H$�QDV�ҡ$��H$�QLVW�ҡ$��H$�AH�U�R�Ћ$��Q�J�E�P�у�_��^��]� �������U��$��P,�E�R@��VWP�E�P�ҋu���$��H�QV�ҡ$��H�QVW�ҡ$��H�A�U�R�Ѓ�_��^��]� ��̡$��H,�j j �҃��������������U��$��P,�EP�EPQ�J�у�]� U��$��H,�AV�u�R�Ѓ��    ^]�������������̡$��P,�B����̡$��P,�B����̡$��P,�B����̡$��P,�B ����̡$��P,�B$����̡$��P,�B(�����U��$��P,�R]�����������������U��$��P,�R��VW�E�P�ҋu���$��H�QV�ҡ$��H$�QDV�ҡ$��H$�QLVW�ҡ$��H$�AH�U�R�Ћ$��Q�J�E�P�у�_��^��]� �������U��$��H��D  ]��������������U��$��H��H  ]��������������U��$��H��L  ]��������������U��$��H�I]�����������������U��$��H�A]�����������������U��$��H�I]�����������������U��$��H�A]�����������������U��$��H�I]�����������������U��$��H���  ]��������������U��$��H�A]�����������������U���V�u�E�P��������$��Q$�J�E�P�у���u-�$��B$�PH�M�Q�ҡ$��H�A�U�R�Ѓ�3�^��]Ë$��Q�J�E�jP�у���u=�U�R��������u-�$��H$�AH�U�R�Ћ$��Q�J�E�P�у�3�^��]Ë$��B�HjV�у���u�$��B�HV�у����I����$��Q$�JH�E�P�ы$��B�P�M�Q�҃��   ^��]�����������U��$��H�A ]�����������������U��$��H�I(]�����������������U��$��H��  ]��������������U��$��H��   ]��������������U��$��H��  ]��������������U��$��H��  ]��������������U��$��H�A$��V�U�WR�Ћ$��Q�u���BV�Ћ$��Q$�BDV�Ћ$��Q$�BLVW�Ћ$��Q$�JH�E�P�ы$��B�P�M�Q�҃�_��^��]������U��$��H���  ��V�U�WR�Ћ$��Q�u���BV�Ћ$��Q$�BDV�Ћ$��Q$�BLVW�Ћ$��Q$�JH�E�P�ы$��B�P�M�Q�҃�_��^��]���U��$��H���  ]��������������U���<�\���SVW�E�    t�E�P�   ��������/�$��Q�J�E�P�   �ы$��B$�PD�M�Q�҃��}�$��H�u�QV�ҡ$��H$�QDV�ҡ$��H$�QLVW�҃���t)�$��H$�AH�U�R����Ћ$��Q�J�E�P�у���t&�$��B$�PH�M�Q�ҡ$��H�A�U�R�Ѓ�_��^[��]���U��$��H�U���  ��VWR�E�P�ы$��u���B�HV�ы$��B$�HDV�ы$��B$�HLVW�ы$��B$�PH�M�Q�ҡ$��H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]���������̡$��H���   ��U��$��H���   V�uV�҃��    ^]�������������U��$��P�]��$��P�B����̡$��P���   ��U��$��P�R`]�����������������U��$��P�Rd]�����������������U��$��P�Rh]�����������������U��$��P�Rl]�����������������U��$��P�Rp]�����������������U��$��P�Rt]�����������������U��$��P���   ]��������������U��$��P�Rx]�����������������U��$��P���   ]��������������U��$��P�R|]�����������������U��$��P���   ]��������������U��$��P���   ]��������������U��$��P���   ]��������������U��$��P���   ]��������������U��$��P���   ]��������������U��$��P���   ]��������������U��$��P���   ]��������������U��$��P���   ]��������������U��$��P���   ]��������������U��$��P���   ]��������������U��$��P�EPQ��  �у�]� �U��$��P���   ]��������������U��$��P���   ]��������������U��$��P���   ]��������������U��E��t �$��R P�B$Q�Ѓ���t	�   ]� 3�]� U��$��P �E�RLQ�MPQ�҃�]� U��E��u]� �$��R P�B(Q�Ѓ��   ]� ������U��$��P�R]�����������������U��$��P�R]�����������������U��$��P�R]�����������������U��$��P�R]�����������������U��$��P�R]�����������������U��$��P�R]�����������������U��$��P�E�R\P�EP��]� ����U��$��E�P�B ���$��]� ���U��$��E�P�B$Q�$��]� �����U��$��E�P�B(���$��]� ���U��$��P�R,]�����������������U��$��P�R0]�����������������U��$��P�R4]�����������������U��$��P�R8]�����������������U��$��P�R<]�����������������U��$��P�R@]�����������������U��$��P�RD]�����������������U��$��P�RH]�����������������U��$��P�RL]�����������������U��$��P�RP]�����������������U��$��P���   ]��������������U��$��P�RT]�����������������U��$��P�EPQ��  �у�]� �U��$��P���   ]��������������U��$��P���   ]��������������U��$��P�RX]����������������̡$��P���   ��U��$��P���   ]��������������U��$��P���   ]��������������U��$��P���   ]��������������U��$��P���   ]�������������̡$��P���   ��U��$��P���   ]�������������̡$��P���   ��$��P���   ��$��P���   ��U��$��H���   ]��������������U��$��H��   ]��������������U��$��H�U�E��VWRP���  �U�R�Ћ$��Q�u���BV�Ћ$��Q�BVW�Ћ$��Q�J�E�P�у�_��^��]������������U��$��H���  ]��������������U��$��P(�BPVW�}�Q�]���E�$�Ѕ�tM�$��G�Q(�]�E�BPQ���$�Ѕ�t,�$��G�Q(�]�E�BPQ���$�Ѕ�t_�   ^]� _3�^]� ����U��$��P(�BTVW�}����$���Ѕ�tE�$��G�Q(�BT�����$�Ѕ�t(�$��G�Q(�BT�����$�Ѕ�t_�   ^]� _3�^]� U��VW�}W��� �����t8�GP���������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U��VW�}W��� �����t8�GP��������t)�O0Q��������t��HW���������t_�   ^]� _3�^]� ������������U��$��} �P(�R8��P��]� ����U��$��P�BdS�]VW��j ���Ћ$��Q�����   hh���h�  V�Ћ$������Eu�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћ$��Q(�BHV���Ѕ�t �$��Q(�E�R VP���҅�t�   �3��EP�`e����_��^[]� ����U���V�E���MP�K���P���#����$��Q�J���E�P�у���^��]� ���U��$��P8�EPQ�JD�у�]� ���̡$��H8�Q<�����U��$��H8�A@V�u�R�Ѓ��    ^]�������������̡$��H8�������U��$��H8�AV�u�R�Ѓ��    ^]��������������U��$��P8�EP�EP�EPQ�J�у�]� ������������U��$��P8�EP�EPQ�J�у�]� �$��P8�BQ�Ѓ����������������U��$��P8�EPQ�J �у�]� ����U��$��P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U��$��P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U��$��P8�EP�EPQ�J(�у�]� U��$��P8�EP�EP�EPQ�J,�у�]� ������������U��$��P8�EP�EP�EPQ�J�у�]� ������������U��$��P8�EP�EP�EP�EP�EPQ�J�у�]� ����U��$��P8�EP�EPQ�J0�у�]� U��$��P8�EP�EP�EPQ�J4�у�]� ������������U��$��P8�EPQ�J8�у�]� ����U��$��H��x  ]��������������U��$��H��|  ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H�A,]�����������������U��$��H�QV�uV�ҡ$��H�Q8V�҃���^]�����̡$��H�Q<�����U��$��H�I@]����������������̡$��H�QD����̡$��H�QH�����U��$��H�AL]�����������������U��$��H�IP]�����������������U��$��H��<  ]��������������U��$��H��,  ]��������������U��$��H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡$��H���   ��$��H���  ��U��$��H�U�ER�UP�ER�UP���   Rh�.  �Ѓ�]����������������U��$��H�A]�����������������U��$��H��\  ]��������������U��$��H�AT]�����������������U��$��H�AX]�����������������U��$��H�A\]����������������̡$��H�Q`����̡$��H�Qd����̡$��H�Qh�����U��$��H�Al]�����������������U��$��H�Ap]�����������������U��$��H�At]�����������������U��$��H��D  ]��������������U��$��H��  ]��������������U��$��H�Ix]�����������������U��$��H��@  ]��������������U��V�u�������$��H�U�A|VR�Ѓ���^]���������U��$��H���   ]��������������U��$��H��h  ]��������������U��$��H��d  ]��������������U��$��H���  ]�������������̡$��H���   ��U��$��H��l  ]��������������U��$��H��   ]��������������U��$��H��  ]��������������U��V�u���R  �$��H���   V�҃���^]���������̡$��H��`  ��U��$��H��  ]��������������U��$��H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U��$��H���  ]��������������U��U�E�$��H�E���   R���\$�E�$P�у�]�U��$��H���   ]��������������U��$��H���   ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H���   ]��������������U��$��H���   ]��������������U��$��H���   ]��������������U��$��H���   ]��������������U��$��H���   ]��������������U��$��H���   ]��������������U��$��P���E�P�E�P�E�PQ���   �у����#E���]����������������U��$��P���E�P�E�P�E�PQ���   �у����#E���]����������������U��$��P���E�P�E�P�E�PQ���   �у����#E���]����������������U��$��H��8  ]��������������U��V�u(V�u$�E�@�$��R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@�$��R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��$��P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U��$��P0�EP�EP�EP�EPQ���   �у�]� ����̡$��P0���   Q�Ѓ�������������U��$��P0�EP�EPQ���   �у�]� �������������U��$��P0�EP�EP�EP�EPQ���   �у�]� ����̡$��P0���   Q�Ѓ������������̡$��H0���   ��U��$��H0���   V�u�R�Ѓ��    ^]�����������U��$��H��H  ]��������������U��$��H��T  ]�������������̡$��H��p  ��$��H���  ��U��$��H���  ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H�U�E��X  ��VR�UPR�E�P�ыu�    �F    �$����   �Qj PV�ҡ$����   ��U�R�Ѓ� ��^��]��������U���$Vj hLGOg�M���  P�E�hicMCP�k������M���  �$����   �JT�E�P�у���u(�u���j  �$����   ��M�Q�҃���^��]á$����   �AT�U�R�Ћu��P���j  �$����   �
�E�P�у���^��]�������������U��$��H��  ]��������������U��$��H��\  ]��������������U��$��H�U��t  ��V�uVR�E�P�у����s����M�������^��]�����U��$��H�U���  ��VWR�E�P�ы$��u���B�HV�ы$��B�HVW�ы$��B�P�M�Q�҃�_��^��]����������������U��$��H�U���  ��VWR�E�P�ы$��u���B�HV�ы$��B�HVW�ы$��B�P�M�Q�҃�_��^��]����������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H�U�E��VWj R�UP�ERP��t  �U�R�Ћ$��Q�u���BV�Ћ$��Q�BVW�Ћ$��Q�J�E�P�у�(_��^��]��U��$��H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    �$����   j P�BV�Ћ$����   �
�E�P�у�$��^��]���U��$��H��8  ]��������������U���  �`�3ŉE��M�EPQ������h   R���  ����|	=�  |#��$��H��0  h��hF  �҃��E� �$��H��4  ������RhЕ�ЋM�3̓�蕉  ��]�������U��$��H��  ��V�U�WR�Ћ$��Q�u���BV�Ћ$��Q�BVW�Ћ$��Q�J�E�P�у�_��^��]����U��$��H��  ��V�U�WR�Ћ$��Q�u���BV�Ћ$��Q�BVW�Ћ$��Q�J�E�P�у�_��^��]����U��$��H��p  ��$�҅�trh���M��  �$��P�E�R4Ph���M��ҡ$��P�E�R4Ph���M���j �E�P�M�hicMCQ�����$����   ��M�Q�҃��M��  ��]�U��$��H��p  ��$V�҅�u�$��H�u�QV�҃���^��]�Wh!���M���
  �$��P�E�R4Ph!���M���j �E�P�M�hicMCQ�����$����   �QHP�ҋu���$��H�QV�ҡ$��H�QVW�ҡ$����   ��U�R�Ѓ�$�M��
  _��^��]������U��$��H��p  ��$V�҅�u�$��H�u�QV�҃���^��]�Wh����M��,
  �$��P�E�R4Ph����M���j �E�P�M�hicMCQ�����$����   �QHP�ҋu���$��H�QV�ҡ$��H�QVW�ҡ$����   ��U�R�Ѓ�$�M���	  _��^��]������U��$��H��p  ��$�҅�u��]�Vh#���M��t	  �$��P�E�R4Ph#���M���j �E�P�M�hicMCQ������$����   �Q8P�ҋ�$����   ��U�R�Ѓ��M��U	  ��^��]���������������U��$��H��p  ��$�҅�u��]�Vhs���M���  �$��P�E�R4Phs���M���j �E�P�M�hicMCQ�W����$����   �Q8P�ҋ�$����   ��U�R�Ѓ��M��  ��^��]���������������U��$��H���  ]��������������U��$��H��@  ]��������������U��$��H���  ]��������������U��V�u���t�$��QP��D  �Ѓ��    ^]������U��$��H��H  ]��������������U��$��H��L  ]��������������U��$��H��P  ]��������������U��$��H��T  ]��������������U��$��H��X  ]��������������U��$��H��\  ]�������������̡$��H��d  ��U��$��H��h  ]��������������U��$��H��l  ]�������������̡$��H���  ��U��$��H�U���  ��VR�E�P�ыu��P���  �M��  ��^��]�����U��$��H���  ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H���  ]��������������U��$��H��$  ]��������������U��$��H��(  ]��������������U��$��H��,  ]�������������̡$��H��0  ��$��H��<  ��U��$��H���  ]�������������̡$��H���  ��U��$��H���  ]������������������������������U��$��H��  ]�������������̡$��H��P  ��$����   ���   ��Q��Y��������U��$��H�A�U��� R�Ћ$��Q�Jj j��E�hԕP�ыUR�E�P�M�Q�m���$��B�P�M�Q�ҡ$��H�A�U�R�Ћ$��Q�J�E�P�у�,��]�̡$��H\�������U��$��H\�AV�u�R�Ѓ��    ^]�������������̡$��P\�BQ�Ѓ���������������̡$��P\�BQ�Ѓ����������������U��$��P\�EPQ�J�у�]� ����U��$��P\�EP�EPQ�J�у�]� U��$��P\�EPQ�J�у�]� ���̡$��P\�BQ�Ѓ����������������U��$��P\�EPQ�J �у�]� ����U��$��P\�EP�EPQ�J$�у�]� U��$��P\�EP�EP�EPQ�J(�у�]� ������������U��$��P\�EPQ�J0�у�]� ����U��$��P\�EPQ�J@�у�]� ����U��$��P\�EPQ�JD�у�]� ����U��$��P\�EPQ�JH�у�]� ���̡$��P\�B4Q�Ѓ����������������U��$��P\�EP�EPQ�J8�у�]� U��$��P\�EPQ�J<�у�]� ����U���SVW�}��j �ωu������$��H\�QV�҃���S������3���~?��I �$��H\�U�R�U��EP�A(VR�ЋM��Q���X����U�R���M�����;�|�_^[��]� �������������U���VW�}�E��P�������}� ��   �$��Q\�BV�Ѓ��M�Q���q����E���taS3ۅ�~L�I �UR���U����E�P���J����E;E�#���$��Q\P�BV�ЋE����;E��E~߃�;]�|�[_�   ^��]� _�   ^��]� �����������̡$��P�BVj j����Ћ�^���������U��$��P�E�RVj P���ҋ�^]� U��$��P�E�RVPj����ҋ�^]� �$��P�B�����U��$��P���   Vj ��Mj V�Ћ�^]� �����������U��$��P�EPQ�J�у�]� ����U��$��P�EPQ�J�у������]� �������������U��$��P�E�RtP�ҋ$����   P�BX�Ѓ�]� ���U��$��P�E�Rlh#  P�EP��]� ���������������U��$��P�E�RlhF  P�EP��]� ���������������U��$��P�E�RtP�ҋ$����   �M�R`QP�҃�]� ���������������U��$��P���   ]��������������U��$��P�E���   P�҅�u]� �$����   P�B�Ѓ�]� �������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������U���   V���  �����   �ESP�M��X����$��Q�J�E�P�ы$��B�Pj j��M�hДQ�҃��E�P�M�����j j��M�Q�U�R��d���P�������P�M�Q�׿����P�U�R�ʿ�����P�  ���M����Q����M��I�����d����>����M��6����$��H�A�U�R�Ѓ��M�������[t	V��  ����^��]� ���U��EVP���!'  �����^]� �����Q�  Y���������U��E�M�U�H4�M�P �U��M�@�] �@8� �@<�P�@@p� �@DpP�@H@� �@L � �@P�P�@l� �@X�P�@\�P�@`�P�@d�P�@T�� �@hP� �@p�� �@t�P�P0�H(�@,    ]��������������U���   h�   ��`���j P��r  �M�U�Ej Q�MRPQ��`���R�����E �Uh�   ��`���Q�E��ERPj�5�����8��]��������������̋�`����������̋�` ����������̋�`0����������̋�`@����������̋�`4����������̋�`����������̋�`8����������̋�`,�����������hD�PhD �`  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d��������]� ���������U��hD�jhD �  ����t
�@��t]��3�]��������VhD�j\hD ���\  ����t�@\��tV�Ѓ���^�����VhD�j`hD ���,  ����t�@`��tV�Ѓ�^�������U��VhD�jdhD ����  ����t�@d��t
�MQV�Ѓ�^]� ������������U��VhD�jhhD ���  ����t�@h��t
�MQV�Ѓ�^]� ������������VhD�jlhD ���|  ����t�@l��tV�Ѓ�^�������U��VhD�h�   hD ���F  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��VhD�h�   hD ����  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��VhD�jphD ���  ����t�@p��t�MQV�Ѓ�^]� �H�^]� ��U��VhD�jxhD ���i  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��VhD�j|hD ���)  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��VhD�j|hD ����  ����t�@|��t�MVQ�Ѓ������^]� �   ^]� ����������̋���������������hD�jhD �  ����t	�@��t��3��������������U��V�u�> t+hD�jhD �S  ����t�@��tV�Ѓ��    ^]�������U��VW�}����t0hD�jhD �  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��VhD�jhD ����  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��VhD�jhD ���  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����VhD�j hD ���L  ����t�@ ��tV�Ѓ�^�3�^���VhD�j$hD ���  ����t�@$��tV�Ѓ�^�3�^���U��VhD�j(hD ����  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��VhD�j,hD ���  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��VhD�j(hD ���Y  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������VhD�j4hD ���  ����t�@4��tV�Ѓ�^�3�^���U��VhD�j8hD ����  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��VhD�j<hD ���  ����t�@<��t
�MQV�Ѓ�^]� ������������VhD�jDhD ���L  ����t�@D��tV�Ѓ�^�3�^���U��VhD�jHhD ���  ����t�M�PHQV�҃�^]� U��VhD�jLhD ����  ����u^]� �M�PLQV�҃�^]� �����������U��VhD�jPhD ���  ����u^]� �M�U�@PQRV�Ѓ�^]� �������VhD�jThD ���l  ����u^Ë@TV�Ѓ�^���������U��VhD�jXhD ���9  ����t�M�PXQV�҃�^]� U��VhD�h�   hD ���  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��VhD�h�   hD ���
  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��VhD�h�   hD ���f
  ����u^]� �M���   QV�҃�^]� �����U��VhD�h�   hD ���&
  ����u^]� �M���   QV�҃�^]� �����U��VhD�h�   hD ����	  ����u^]� �M���   QV�҃�^]� �����U��VhD�h�   hD ���	  ����t�M�UQ�MR���   QV�҃�^]� ��U���VhD�h�   hD �e	  ����u�$��H�u�QV�҃���^��]ËM���   WQ�U�R�Ћ$��Q�u���BV�Ћ$��Q�BVW�Ћ$��Q�J�E�P�у�_��^��]��U��VhD�h�   hD ����  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��VhD�h�   hD ���  ����t���   ��t�MQ����^]� 3�^]� �U��VhD�h�   hD ���F  ����t���   ��t�MQ����^]� 3�^]� �U��VhD�h�   hD ���  ����t���   ��t�MQ����^]� 3�^]� �VhD�h�   hD ����  ����t���   ��t��^��3�^����������������U��VhD�h�   hD ���  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��VhD�h�   hD ���6  ����t���   ��t�MQ����^]� ��������U��VhD�h�   hD ����  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������VhD�h�   hD ���  ����t���   ��t��^��3�^����������������VW��3����$    �hD�jphD �_  ����t�@p��t	VW�Ѓ���H��8 t����_��^�����U��SW��3�V��    hD�jphD �  ����t�@p��t	WS�Ѓ���H��8 tshD�jphD ��  ����t�@p��t�MWQ�Ѓ�����H�hD�jphD �  ����t�@p��t	WS�Ѓ���H�V���7�����t���[����E��^t�8��~=hD�jphD �\  ����t�@p��t	WS�Ѓ���H��8 u_�   []� _3�[]� ��������U��VhD�j\hD ���	  ����t3�@\��t,V��hD�jxhD ��  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��VhD�j\hD ���  ����t3�@\��t,V��hD�jdhD �  ����t�@d��t
�MQV�Ѓ���^]� ��������U���VhD�j\hD ���F  ����tG�@\��t@V�ЋEhD�jdhD �E��E�    �E�    �  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��VhD�j\hD ����  ����t\�@\��tUV��hD�jdhD �  ����t�@d��t
�MQV�Ѓ�hD�jhhD �~  ����t�@h��t
�URV�Ѓ���^]� ���������������U��VhD�j\hD ���9  ������   �@\��t~V��hD�jdhD �  ����t�@d��t
�MQV�Ѓ�hD�jhhD ��  ����t�@h��t
�URV�Ѓ�hD�jhhD ��  ����t�@h��t
�MQV�Ѓ���^]� ��U���VhD�jthD ���  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���hD�j`hD �N  ����t(�@`��t!�M�Q�Ѓ���^��]� �uhH����_�����^��]� ������U���VhD�h�   hD ����  ����tR���   ��tH�MQ�U�R���ЋuP������hD�j`hD �  ����t<�@`��t5�M�Q�Ѓ���^��]� �u�U�R���E�    �E�    �E�    ������^��]� ��������������U��$����   �BXQ�Ѓ���u]� �$��Q|�M�RQ�MQP�҃�]� ���U��$����   �BXQ�Ѓ���u]� �$��Q|�M�R8Q�MQP�҃�]� ���U��EV��j ��$��Qj j P�B�ЉF����^]� ��̡$�Vj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� �$��Q�MP�EP�Q�JP�у��F�   ^]� ����U��E�M�UP��P�EjP������]��������������̸   �����������U��V�u��t���u8�EjP��������u3�^]Ë��������t���t��U3�;P����#�^]�����U��M�EV�u������t#W���    �Pf�y������f�8f�u�_^]� �U��� �E���M��"  �ȉES���V�u��W�}�ǃ��Q���ƃ��։E��B��E���؉M�E��U���M��~�U�U���)}�M��>���E��}�t�u+���I �\�P���m���u�E�����E��   )}��u��	;]��u��s���u;]�]�}�M��>P�E�V�Ѕ�}	�u���]�M��E��VP�҅��V������F��}�t!�M�+ȃ����\�P���m���u�]��;]~�����_^[��]� ���U���(W�}�����E�E���M��  �MS�؉E������ǃ��S�����E�ы���V�]�U��E܉U���]��~�E�E��)}��]��)�M�U��E�Q�M�RP������E�����E��   )}��u�;E��؉u�s���u;]�]�}�M���>P�E؋V�Ѕ�}	�u؃��]��M���E�VP�҅��i����}���F�t&�M�+ȃ���I �Pf�\����f�f�u�]��}�;E�w����%���^[_��]� ��������U���(W�}�����E�E���M��)  �ЉE������ǃ��J���SV�uƃ��ΉE��A��E����؉U��E܉M����I �U���~�M�M��)}��U��A�M�ɋE��M�t�M�+���I �\�p���m���4u�E�����E��   )}��u�;E��؉u�s���u;]�]�}�M��>P�E؋V�Ѕ�}	�u؃��]��M��E�VP�҅��Q����}���F�t�M�+ȃ���\�P������u�]��}�;E~�����^[_��]� ���������������U��E�Pu�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����E��SV��W�]�t8�u��t1�}��t*�} t$�VP��Ѕ���   |������E�   �}}_^3�[��]� �}�M���E�������uu��VP�҅�t#}����}����}��E9E�~�_^3�[��]� ��~3�E���]��]�E��E�M���؋ESP���҅�u�����_��^[��]� ���������������U����E��SV��W�]��  �u����   �}����   �} ��   �VP��Ѕ���   }�M_^�    3�[��]� �O�3����E�   �M} ����   �E���8_^3�[��]� ���M�U���<�M������uuVQ���҅�t}�O��M��W�U��M9M�~�뤅�~3�E���]��]�E��E�M���؋ESP���҅�u�����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� ����������̡$��H���   ��U��$��H���   V�u�R�Ѓ��    ^]����������̡$��P���   Q�Ѓ�������������U��$��P�EPQ���   �у�]� ̡$��H�������U��$��H�AV�u�R�Ѓ��    ^]��������������U��$��H�AV�u�R�Ѓ��    ^]��������������U��$��P��Vh�  Q���   �E�P�ы$����   �Q8P�ҋ�$����   ��U�R�Ѓ���^��]��������������̡$��P�BQ�Ѓ����������������U��$��P�EPQ�J\�у�]� ����U��$��P�EP�EP�EP�EP�EPQ���   �у�]� �U��$��P�EP�EP�EP�EPQ�JX�у�]� �������̡$��P�B Q��Y�U��$��P�EP�EP�EP�EPQ���   �у�]� �����U��$��P�EP�EP�EPQ�J�у�]� ������������U��$��H��   ]��������������U��$��P�R$]�����������������U��$��P��x  ]��������������U��$��P�EP�EP�EP�EPQ�J(�у�]� ��������U��$��P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U��$��P�EP�EP�EP�EPQ�J,�у�]� ��������U��$�V��H�QWV�ҋ��$��H�QV�ҋ$��Q�M�R4Q�MQ�MQ���W���Pj j V�҃�(_^]� �����������U��$��P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U��$��P�EP�EPQ�J@�у�]� U��$��P�EPQ�JD�у�]� ���̡$��P�BLQ�Ѓ���������������̡$��P�BLQ�Ѓ���������������̡$��P�BPQ�Ѓ����������������U��$��P�EPQ�JT�у�]� ����U��$��P�EPQ�JT�у�]� ����U��$��P�EP�EPQ���   �у�]� �������������U��$��P�E���   ��VP�EPQ�M�Q�ҋu�    �F    �$����   j P�BV�Ћ$����   �
�E�P�у� ��^��]� ������̡$��P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡$��H�������U��$��H�AV�u�R�Ѓ��    ^]��������������U��$��P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U��$��P�EPQ�J�у�]� ���̡$��P�BQ��Y�U��$��P�EP�EPQ�J�у�]� U��VW��������M�U�x@�EPQR�������H ���_^]� �U��VW�������M�U�xD�EPQR���~����H ���_^]� �V���h����xH u3�^�W���V����΍xH�L����H �_^�����U��V���5����xL u3�^]� W��� ����M�U�xL�EPQR���
����H ���_^]� �������������U��V��������xP u���^]� W��������M�U�xP�EP�EQRP�������H ���_^]� ��������U��V�������xT u���^]� W�������M�xT�EPQ���m����H ���_^]� U���S�]��VW��t.�M��V������?����xL�E�P���1����H ��ҍM������}��tZ�$��H�A�U�R�Ћ$��Q�J�E�WP�ы$��B�P�M�Q�҃���������@@��t�$��QWP�B�Ѓ�_^[��]� ������U��V�������x` u
� }  ^]� W�������x`�EP�������H ���_^]� ��U��VW���d����xH�EP���V����H ���_^]� ���������U��SVW���3����x` u� }  �#�������x`�E���P�������H ��ҋ��$��H�]�QS�҃�;�A�$��H�QS�҃�;�,��������M�U�xD�EPQSR�������H ���_^[]� _^�����[]� ��������������U��V�������xP u
�����^]� W���m����M�U�xP�EP�EQ�MR�UPQR���K����H ���_^]� ��������������U��V���%����xT u
�����^]� W�������M�xT�EPQ��������H ���_^]� ��������������U��V��������xX tW��������xX�EP�������H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u��H=  ����t.�E�;�t'�$��J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡$��H��   ��U��$��H��$  V�u�R�Ѓ��    ^]�����������U��$��UV��H��(  VR�Ѓ���^]� �����������U��$��P�EQ��,  P�у�]� �U��$��P�EQ��,  P�у������]� ���������̡$��H��0  ��$��H��4  ��$��H��p  ��$��H��t  ��U��E��t�@�3��$��RP��8  Q�Ѓ�]� �����U��$��P�EPQ��<  �у�]� �U��$��P�EP�EP�EPQ��@  �у�]� ���������U��$��P�EP�EPQ��D  �у�]� �������������U��$��P�EPQ��H  �у�]� �U��$��P�E��L  ��VWPQ�M�Q�ҋu���$��H�QV�ҡ$��H�QVW�ҡ$��H�A�U�R�Ѓ�_��^��]� ��������������̡$��P��T  Q�Ѓ�������������U��$��P�EPQ��l  �у�]� ̡$��P��P  Q�Ѓ�������������U��$��P�EPQ��X  �у�]� ̡$��H��\  ��U��$��H��`  V�u�R�Ѓ��    ^]�����������U��$��P�EP�EP�EP�EP�EPQ��d  �у�]� �U��$��P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���w��������3��F�F �F$�F(�F,�F0�F4�F8�F<�F@�FD�FH�FL�FP�FT�FX�_p��G`�Gd�Gh�Gx�����G|   ��_^��������������V��W�>��t7���O����xP t$S���A���j j �XPj�FP���-����H ���[�    �~` t�$��H�V`�AR�Ѓ��F`    _^������������U��SV��Fx�$��Q��   WV�^dSP�EP�~`W�у����F|��   �> ��   �; ��   �U�~pW�^hSR�Ĺ������u#���hؕ�$��H��0  h�   �҃��E�~P��輒���j j jW�^������F|t��������F|_^[]� �F|_�Fx����^[]� �F|�����    �$��Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��V��~d �F`tLW�};~xtBWPj�NQ��������F|u�E���~xt�    �F`_^]� �M���Fx����t�3�_^]� U��QVW�}����9  �$��H�QhV�҃����$�u"�H��0  hؕh�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���t�3�9u�~!�E���<� t��Q���_7  �E��;u�|�UR�����_�   ^��]� �����������U��QVW�}�����8  �$��H�QhV�҃����$�u"�H��0  hؕh�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���tЋE��t�3�9u�~:��E�<� t'���$��QP�Bh�Ѓ���t�M��R���|6  ��;u�|ȍEP�����_�   ^��]� �����������hؕh�   hp�h�   �������t�������3��������V���(����N^鯌�����������������U��VW�}�7��t��������N背��V�m�����    _^]Ë�3ɉH��H�@   �������������U��ыM��tK�E��t�$����   P�B@��]� �E��t�$����   P�BD��]� �$����   R�PD��]� �����U��$��P@�Rd]�����������������U��$��P@�Rh]�����������������U��$��P@�Rl]�����������������U��$��P@�Rp]�����������������U��$����   ���   ]�����������U��$����   ���   ]����������̡$��P@�Bt����̡$��P@�Bx�����U��$��P@�R|]����������������̡$��P@���   ��$����   �Bt��U��$��P@���   ]�������������̡$��P@���   ��U��$��P@���   ]��������������U��$��P@���   ]��������������U��$��P@���   ]��������������U��$��P@���   ]��������������U��$�V��H@�QV�ҋM����t��#����$��Q@P�BV�Ѓ�^]� �̡$��PH���   Q�Ѓ�������������U��$��P@�EPQ�JL�у�]� ���̡$��P@�BHQ�Ѓ����������������U��$��P@�EP�EP�EPQ�J�у�]� ������������U��$��P@�EPQ�J�у�]� ����U��$��P@�EP�EPQ�J�у�]� U��$��P@�EPQ�J �у�]� ����U��$����   �R]��������������U��$����   �R]��������������U��$����   �R ]��������������U��$����   ���   ]�����������U��$����   ��D  ]�����������U��$��E���   �E ���   P�E���$P�EP�EP�EP��]� ���������U��$����   ���   ]����������̡$����   �B$��$��H@�Q0�����U��$��H@�A4j�URj �Ѓ�]����U��$��H@�A4j�URh   @�Ѓ�]�U��$��H@�U�E�I4RPj �у�]�̡$��H|�������U��V�u���t�$��Q|P�B�Ѓ��    ^]��������̡$��H|�Q �����U��V�u���t�$��Q|P�B(�Ѓ��    ^]��������̡$��H@�Q0�����U��V�u���t�$��Q@P�B�Ѓ��    ^]���������U��$��H@���   ]��������������U��V�u���t�$��Q@P�B�Ѓ��    ^]��������̡$��PH���   Q�Ѓ�������������U��$��PH�EPQ��d  �у�]� �U��$��H �IH]�����������������U��}qF uHV�u��t?�$����   �BDW�}W���Ћ$��Q@�B,W�Ћ$��Q�M�Rp��VQ����_^]����������̡$��P@�BT�����U��$��P@�RX]�����������������U��$��P@�R\]����������������̡$��P@�B`�����U��$��H��T  ]��������������U��$��H@�U�A,SVWR�Ћ$��Q@�J,���EP�ы$��Z��h��hE  �΋��6���Ph��hE  ���$���P��T  �Ѓ�_^[]����hT�Ph^� ��������������������U��VhT�jh^� ����������t�@��t�M�UQRV�Ѓ�^]� 3�^]� �VhT�jh^� ���|�������t�@��tV�Ѓ�^�3�^���U��VhT�jh^� ���I�������t�@��t�M�UQRV�Ѓ�^]� ���^]� U���  VhT�jh^� ����������t/�@��t(�MWQ��x���VR�Ћ��E���b   ���_^��]� �u�������N`�������   ������   ������ݞ�  ��^��]� ����U��VhT�jh^� ���y�������t�@��t�M�UQRV�Ѓ�^]� ��������U��VhT�jh^� ���9�������t�@��t�M�UQ�MRQV�Ѓ�^]� ����U��VhT�j h^� �����������t�@ ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��VhT�j$h^� ����������t�@$��t�MQV�Ѓ�^]� 3�^]� �����U��VhT�j(h^� ���i�������t�@(��t�M�UQ�MR�UQRV�Ѓ�^]� U��QVhT�j,h^� ���(�������t �@,���E�t�E�MPQV�U���^��]� ��^��]� ��������U��VhT�j0h^� �����������t#�@0��t�E�M�U���$QRV�Ѓ�^]� 3�^]� ��������VhT�j4h^� ����������t�@4��tV�Ѓ�^�3�^���VhT�j8h^� ���\�������t�@8��tV�Ѓ�^�������U���`VhT�jDh^� ���&�������t(�@D��t!W�M�VQ�Ћ��E���   ���_^��]� �u�������^��]� ����U��VhT�jHh^� �����������t�@H��t
�MQV�Ѓ�^]� ������������U��VhT�jLh^� ����������t�@L��t�MQV�Ѓ�^]� ���^]� ����U��VhT�jPh^� ���I�������t�@P��t
�MQV�Ѓ�^]� ������������U��VhT�jTh^� ���	�������t�@T��t
�MQV�Ѓ�^]� ������������U��VhT�jXh^� �����������t.�@X��t'�M �UQ�MR�UQ�MR�UQ�MRQV�Ѓ� ^]� 3�^]� �������������VhT�j`h^� ���l�������t�@`��tV�Ѓ�^�3�^���U��VhT�jdh^� ���9�������t�@d��t�MQV�Ѓ�^]� 3�^]� �����U���VhT�jhh^� �����������t1�@h��t*�MQ�U�VR�Ћu��P�������M�������^��]� �u���D�����^��]� �����������VhT�jph^� ����������t�@p��tV�Ѓ�^Ã��^��VhT�jlh^� ���\�������t�@l��tV�Ѓ�^Ã��^��VhT�jth^� ���,�������t�@t��tV�Ѓ�^�3�^���U��VhT�jxh^� �����������t�@x��t
�MQV�Ѓ�^]� ������������VhT�j|h^� ����������t�@|��tV�Ѓ�^�������VhT�h�   h^� ����������t���   ��tV�Ѓ�^�U��VhT�h�   h^� ���V�������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������U��VhT�h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U���VhT�h�   h^� ����������tU���   ��tKW�M�VQ�Ћ$��u���B�HV�ы$��B�HVW�ы$��B�P�M�Q�҃�_��^��]� �$��H�u�QV�҃���^��]� ����������VhT�h�   h^� ����������t���   ��tV�Ѓ�^Ã��^������������U��VhT�h�   h^� �����������t���   ��t
�MQV�Ѓ�^]� ������U��VhT�h�   h^� ����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��VhT�h�   h^� ���F�������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������VhT�h�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������U��VhT�h�   h^� ����������t%���   ��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���U��VhT�h�   h^� ���f�������t���   ��t�M�UQRV�Ѓ�^]� ���^]� ����������U��VhT�h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��VhT�h�   h^� �����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��VhT�h�   h^� ���v�������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��VhT�h�   h^� ���&�������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������VhT�h�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������VhT�h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������VhT�h�   h^� ���Y�������t���   ��tV�Ѓ�^�3�^�������������VhT�h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������U��VhT�h�   h^� �����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������VhT�h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������U���VhT�h�   h^� ���C�������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��VhT�h�   h^� �����������t���   ��t�M�UQRV�Ѓ�^]� ��VhT�h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������U���VhT�h�   h^� ���C�������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��VhT�h�   h^� �����������t���   ��t�M�UQRV�Ѓ�^]� ��VhT�h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������U��VhT�h�   h^� ���F�������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��QVhT�h�   h^� �����������t#���   ���E�t�E�MPQV�U���^��]� ��^��]� ��U��VhT�h�   h^� ����������t!���   ��t�E�M�U���$QRV�Ѓ�^]� ���������U��VhT�h�   h^� ���V�������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��VhT�h�   h^� ����������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��VhT�h   h^� ����������t��   ��t�MQV�Ѓ�^]� 3�^]� ���������������VhT�h  h^� ���i�������t��  ��tV�Ѓ�^�3�^�������������U���VhT�h  h^� ���#�������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���VhT�h  h^� ����������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���VhT�h  h^� ���#�������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U��VhT�h  h^� ����������t��  ��t
�MQV�Ѓ�^]� ������U��VhT�h  h^� ���f�������t��  ��t
�MQV�Ѓ�^]� ������U��VhT�h  h^� ���&�������t��  ��t
�MQV�Ѓ�^]� ������VhT�h   h^� �����������t��   ��tV�Ѓ�^�3�^�������������U��VhT�h$  h^� ����������t��$  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��VhT�h(  h^� ���V�������t!��(  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��VhT�h,  h^� ����������t��,  ��t�M�UQ�MRQV�Ѓ�^]� ��������������VhT�h0  h^� ����������t��0  ��tV�Ѓ�^�3�^�������������U��VhT�h4  h^� ���v�������t��4  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��VhT�h8  h^� ���&�������t��8  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��VhT�h<  h^� �����������t��<  ��t�M�UQ�MRQV�Ѓ�^]� ��������������U��VhT�h@  h^� ����������t��@  ��t�M�UQ�MRQV�Ѓ�^]� ��������������VhT�hD  h^� ���9�������t��D  ��tV�Ѓ�^�3�^�������������U��VhT�hH  h^� �����������t��H  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��VhT�hL  h^� ����������t��L  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��VhT�hP  h^� ���V�������t!��P  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��QVhT�hT  h^� ����������t'��T  ���E�t�E�M�UPQRV�U���^��]� ��^��]� ��������������U��VhT�hX  h^� ����������t%��X  ��t�E�M�U���$Q�MRQV�Ѓ�^]� �����U��VhT�j<h^� ���Y�������t�@<��t�M�UQRV�Ѓ�^]� ��������U��VhT�j@h^� ����������t�@@��t�MQV�Ѓ�^]� 3�^]� �����hX�Ph�� ��������������������hX�jh�� ��������uË@����U��V�u�> t/hX�jh�� ��������t��U�M�@R�Ѓ��    ^]���U��VhX�jh�� ���Y�������t �@��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��VhX�jh�� ���	�������t�@��t�M�UQR����^]� ����������U��VhX�jh�� �����������t�@��t�M�UQR����^]� ����������U��VhX�jh�� ����������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��VhX�j h�� ���9�������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��VhX�j$h�� �����������t �@$��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��VhX�j(h�� ����������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��VhX�j,h�� ���I�������t0�@,��t)�M$�E�UQ�M���\$�E�$R�UQR����^]�  3�^]�  �����������U��VhX�j0h�� �����������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��VhX�j4h�� ����������t5�@4��t.�M(�E �UQ�M���$R�UQ�MR�UQ�MRQ����^]�$ 3�^]�$ ������U��QVhX�j8h�� ���8�������t�@8���E�t�E�MPQ���U�^��]� ��^��]� ����������U��VhX�j<h�� �����������t�@<��t�M�UQR����^]� ����������U��VhX�j@h�� ����������t�@@��t�M�UQR����^]� 3�^]� ���U��VhX�jHh�� ���i�������t�@H��t�M�UQR����^]� 3�^]� ���U��VhX�jDh�� ���)�������t�@D��t�M�UQR����^]� 3�^]� ���U��QVhX�jLh�� ����������t#�@L���E�t�E�EP�����$�U�^��]� ��^��]� �����U��VhX�jPh�� ��虿������t�@P��t�M�UQR����^]� 3�^]� ���U��VhX�jTh�� ���Y�������t �@T��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��VhX�jXh�� ���	�������t(�@X��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��VhX�j\h�� ��蹾������t(�@\��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��V��~ Wu hX�jh�� �b�������t�@�ЉF�~��t6hX�jh�� �;�������t�@��t�M�UVQ�MRQ����_^]� _3�^]� ��������������U��V��W�~��t+hX�jh�� ��������t�@��t�M�UQR���Ѓ~ t1hX�jh�� 谽������t�N�U�M�@R�Ѓ��F    _^]� ����������U��V��~ u hX�jh�� �c�������t�@�ЉF�v��t+hX�jh�� �<�������t�@��t�M�UQR����^]� �������������U��V�q��t@hX�jh�� ���������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ��������������U��V�q��t<hX�j h�� 蔼������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U��SV��~ Wu hX�jh�� �A�������t�@�ЉF�}�]�M�UWSQR���[�����t�N��t�E�UWSPR����_^[]� _^3�[]� �U��V�q��t8hX�j(h�� �Ի������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� ������U��I��t)�E$�E�UP�E���\$�E�$R�UPR����]�  3�]�  �������U��V�q��t<hX�j0h�� �D�������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �̡$��PD�BQ�Ѓ���������������̡$��PD�BQ�Ѓ���������������̡$��PD�BQ�Ѓ����������������U��$��PX��Q�
�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ���������U��$��PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U��$��PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U��$��PX��`VWQ�J�E�P�ы��E���   ���_^��]� �������������U��$��PX�EPQ�J�у�]� ����U��$��PX�EPQ�J�у�]� ����U��$��PX�EPQ�J�у�]� ����U��$��PX�EPQ�J�у�]� ����U��$��PX�EPQ�J$�у�]� ����U��$��PX�EPQ�J �у�]� ����U��$��PD�EP�EPQ�J�у�]� U��$��HD�U�j R�Ѓ�]�������U��$��H@�AV�u�R�Ѓ��    ^]��������������U��$��HD�	]��U��$��H@�AV�u�R�Ѓ��    ^]��������������U��$��HD�U�j R�Ѓ�]�������U��$��H@�AV�u�R�Ѓ��    ^]��������������U��$��U�HD�Rh2  �Ѓ�]����U��$��H@�AV�u�R�Ѓ��    ^]��������������U��$��U�HD�RhO  �Ѓ�]����U��$��H@�AV�u�R�Ѓ��    ^]��������������U��$��U�HD�Rh'  �Ѓ�]����U��$��H@�AV�u�R�Ѓ��    ^]�������������̡$��HD�j h�  �҃�����������U��$��H@�AV�u�R�Ѓ��    ^]�������������̡$��HD�j h:  �҃�����������U��$��H@�AV�u�R�Ѓ��    ^]��������������U���3��E��E��$����   �R�E�Pj�����#E���]�̡$��HD�j h�F �҃�����������U��$��H@�AV�u�R�Ѓ��    ^]�������������̡$��HD�j h�_ �҃�����������U��$��H@�AV�u�R�Ѓ��    ^]��������������U��E����u��]� �E��$��E�    ���   �R�E�Pj������؋�]� ̡$��PD�B$Q�Ѓ���������������̡$��PD�B(Q�Ѓ���������������̡$��PD�BQ�Ѓ���������������̡$��PD�B(Q�Ѓ���������������̡$��PD�BQ�Ѓ���������������̡$��PD�B(Q�Ѓ���������������̡$��PD�BQ�Ѓ���������������̡$��PD�B(Q�Ѓ���������������̡$��PD�BQ�Ѓ���������������̡$��PD�B(Q�Ѓ���������������̡$��PD�BQ�Ѓ���������������̡$��PD�B(Q�Ѓ���������������̡$��PD�BQ�Ѓ���������������̡$��PD�B(Q�Ѓ���������������̡$��PD�BQ�Ѓ���������������̡$��PD�B(Q�Ѓ���������������̡$��PD�BQ�Ѓ���������������̡$��PD�B(Q�Ѓ���������������̡$��PD�BQ�Ѓ����������������U��E��u�E�M�d��`��   ]� �����������U��E�����V��   �$�ܲ�   ^]áh������h�uT�EP裫����=�.  }�����^]Ëu��t�h�jmhp�j��������t ����W�����\�tV����[���   ^]��\�    �   ^]ËM�UQR��������������^]�^]�����-h�u.�̪��������\���t���fX��V�P������\�    �   ^]Ã��^]Ð������ղr�������������hl�Ph�f �P������������������U��hl�jh�f �,�������t
�@��t]�����]�������U��Vhl�jh�f �����������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R�JW���E�NP�у�4�M���tW����^]ÍM�gW�����^]��U��hl�jh�f 茰������t
�@��t]��3�]��������U��hl�jh�f �\�������t�x t�P]��3�]������V��F��Wu�~��N�ɍ<u�< ��u_3�^á$��H�F��  hL�j8��    RP�у���tщ~�F_�   ^���U��V��F;Fu������u^]� �N�V�E���   F^]� �����������U��V��FW�};�~ ��|�F�M��_�   ^]� _3�^]� })�V;Vu��������t�F�N��    �F9~|׋V;Vu���������t��F�N�U���F_�   ^]� ������U��V��FW�};�~����}3�;Fu������u_^]� �F;�~�N�T������;ǉ�F�M���F_�   ^]� �U��E��|4�Q;�}-���;Q}V�d$ �Q�t������2;A|�^�   ]� 3�]� ������������U��Q3���V~�I�u91t����;�|���^]� �������V��W�~W����3����_�F�F^�����A    ��������̋Q�B���|;�}�QV�4���tP�1�����^�3�����������̍Q3��Q�Q�A�Q�A������������W���O�G;�t#��tV�q��t�~ u3���j�҅���u�^�G�G�G�G    �G�G    _�����U��A��3�;�Vt!��t�M���;�t�@��t
�x t��u�3�^]� ��������U��Q�E�P�Q�P�Q�B�A]� �U��E�Q�P�Q�P�Q�B�A]� ̋Q��3�;�t�ʅ�t�I����t
�y t��u�����������U��E�P�Q�H�A�@�H]� ����U��E�P�Q�H�A�A�H]� ���̋Q��t!�A��t�B�A�Q�P�A    �A    ��������V��W�~W�������3����_�F�F^��������������U���SV�uW���^S�}��f���3���F�F�O�N�W���V9G�E~��I �O���F9F�U�uL��u�~��~��t���< ��t\�$��H���  hL�j8��    RP�у���t3�~�}���V��M����E�F��;G�E|�_^�   [��]� _^3�[��]� �������������U��V�u��|'�A;�} �U��|;�};�t�A��W�<��<���_^]� ���������U��EV�u;�}����|,�Q;�}%��|!;�};�t�QW�<�P������tVW����_^]� ����������U��V�q3���W~�Q�}9:t����;�|���P�����_^]� ���������������U����E�Qj�E��ARP�M��E���諮����]� �����U����Q�Ej�E��A�MRPQ�M��E����Ǯ����]� ̋A��;�t?W3�;�t7V�H;�t	9yt���3��P;�t;�t�J�H�P�Q�x�x;���u�^_������̋Q���H�t!�A��t�B�A�Q�P�A    �A    �̋�� ���@H��HV3��q�q�P�r�r�H��p�p�p�P�H^������V����������F3�;��FH�t�N;�t�H�F�N�H�V�V�F;��FH�t�N;�t�H�F�N�H�V�V^�U��E�UP�AR�Ѓ�]� ���������U��V��N3�;��H�t�F;�t�A�F�N�H�V�V�Et	V�6�������^]� ������������U��V��W�~W��������3����E��F�Ft	V�������_��^]� ������U��V��������Et	V���������^]� ø9��h��l�5��p����t�'��x����|��������������������������"  �|$ �x�t�  ��Ã��$��  �   ��ÍT$�  R��<$�D$tQf�<$t�P  �   �u���=t� ��  �   �0���  �  �u,��� u%�|$ u���%  �"��� u�|$ u�%   �t����-���   �=t� �f  �   �0��o  Z�Q����6  Y�V��������D$tV�c���Y��^� U��Q�E��SVW�  ����   Wj ��P������u3��  V�>����Vj u��P���ދF�~�E�F�E�F�E����  ��P���E��t�� �  �M�����E�����j����������=����.  ��Y�s����!  ��u
�/  �`����
.  ������,  �����&  ��}�t  ����+  ��| �v)  ��|j �$  ��Yu�|��   �
)  ��3�;�u59=|�������|�9=�u�a%  9}u{��(  �  �y.  �j��uY��  h  j��%  ��;�YY�����V�5���5���*  Y�Ѕ�tWV�  YY� ��N���V��  Y�m�����uW�J   Y3�@_^[�� jh����/  ����]3�@�E��u9|���   �e� ;�t��u.�����tWVS�ЉE�}� ��   WVS������E����   WVS�����E��u$��u WPS����Wj S���������tWj S�Ѕ�t��u&WVS�~�����u!E�}� t�����tWVS�ЉE��E������E���E��	PQ��.  YYËe��E�����3��C/  Ã|$u��0  �t$�L$�T$�����Y� QSUVW�5���  �5����t$�  ��;�YY��   ��+ލk��rxV�'1  ��;�YsJ�   ;�s���;�rP�t$�B$  ��YYu�F;�rCP�t$�+$  ��YYt3��P�<���  Y���t$��  ���W�  Y���D$Y�3�_^][Y�Vjj �#  ��V�  ��������ujX^Ã& 3�^�jhе��-  �   �e� �u�����Y�E��E������	   �E��.  ��d   ��t$���������YH�jh��-  �e� �u;5Xw"j�'2  Y�e� V�i:  Y�E��E������	   �E��-  �j�$1  Y�U�l$�����   S��VW3�95$���u�
  j�c  h�   �  YY�l��u;�t���3�@P���uU�S���;�Yu;�u3�G�����WV�5$��Ӌ���u&9��j_tU�"=  ��Yu����<  �8��<  �8_��^[]�U� =  Y�<  �    3�]����̋T$�L$��ti3��D$��u��   r�=L t�9=  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�jh��
,  �u��tu�=luCj�0  Y�e� V�1  Y�E��t	VP� 1  YY�E������   �}� u7�u�
j�/  Y�Vj �5$�����u�;  ����P�d;  �Y��+  ���������U��WV�u�M�}�����;�v;���  ��   r�=L tWV����;�^_u^_]�8=  ��   u������r*��$�t���Ǻ   ��r����$����$�����$���������#ъ��F�G�F���G������r���$�t��I #ъ��F���G������r���$�t��#ъ���������r���$�t��I k�X�P�H�@�8�0�(��D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�t������������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�������$����I �Ǻ   ��r��+��$���$���$�H�p��F#шG��������r�����$���I �F#шG�F���G������r�����$����F#шG�F�G�F���G�������V�������$���I ����������������D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$���� �(�8�L��E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̃=L t-U�������$�,$�Ã=L t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$��;`�u���;  �D$��V���F uc�U  �F�Hl��Hh�N�;�t�$��Hpu�TE  ��F;(�t�F�$��Hpu��=  �F�F�@pu�Hp�F�
���@�F��^� U���V�u�M��l����u�P�H  ��e�F�P��F  ��Yu��P�H  ��xYuFF�M����   �	��	�F�����F��u�8M�^t�E��`p���U���V�u�M�������E��ɋu�t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B�Ɉu��}� ^t�E��`p�����D$�����Az3�@�3��U��QQ�} �u�ut�E�P�CG  �M��E��M��H��EP��G  �E�M�����j �t$�t$�t$������Å�V��tV�K  @PV�V�>H  ��^�j �t$�z���YY�j �t$�����YY�U���SVW�u�M��������3�;�u+�*5  j_VVVVV�8��D  ���}� t�E��`p����!  9uv�9u~�E�3���	9Ew	��4  j"뺀} t�U3�9u��3Ƀ:-����ˋ��:����}�?-��u�-�s�} ~�F�����E����   � � �3�8E��E��}�u����+�]h��SV�4K  ��3ۅ�tSSSSS� C  ��9]�Nt�E�GF�80t.�GHy���-F��d|
�jd_�� ��F��
|
�j
_�� �� F���t�90uj�APQ��F  ���}� t�E��`p�3�_^[��U���,�`�3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�YL  3ۃ�;�u�3  SSSSS�0�=C  �����o�E;�v����uu����3Ƀ}�-��+�3�;���+��M�Q�NQP3��}�-��3�;�����Q�uJ  ��;�t���u�E�SP�u��V�u��������M�_^3�[������U��j �u�u�u�u�u������]�U���$VW�u�M��E��  3��E�0   �k���9}}�}�u;�u+�2  j^WWWWW�0�TB  ���}� t�E�`p����  9}vЋE��9E� w	�}2  j"���}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW� �������t�}� � ��  �M�ap��  �;-u�-F�0F�} je����$�x�FV�6  ��YY�L  �} ���ɀ����p��@ �2  %   �3��t�-F�]�0F������$�x��OF��ۃ����  �3���'3��u!�0�O����� F�u�U���E��  ��1F��F9U�Eu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~M�W#U���M�#E���� �%K  f0 ��f=9 vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� ��J  f= v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V�������u�E�8 u���} �4����$�p���WF�]J  3�%�  #�+E�SY�x;�r�+F�
�-F�����;Ӌ��0|$��  ;�rSQRP�8I  0�F;��U�����u��|��drj jdRP�I  0��U�F����;�u��|��
rj j
RP��H  0��U�F���]�0��F �}� t�E�`p�3�[_^��U���SVW�u�؋s���M�N������u-�\/  j^�03�PPPPP��>  ���}� t�E��`p����   �} v̀} t;uu3��;-����� 0�@ �;-��u�-�w�C3�G�����n����0F���} ~D���Y����E����   � � ��[F��}&�ۀ} u9]|�]�}���(���Wj0V�������}� t�E��`p�3�_^[��U���,�`�3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�G  3ۃ�;�u�O.  SSSSS�0��=  �����Z�E;�v���u��3Ƀ}�-��+��u�M�Q�M��QP3��}�-���P�4E  ��;�t���u�E�SV�u���d������M�_^3�[�b�����U���0�`�3ŉE��ESV�uWj_W�M�Q�M�Q�p�0�NF  3ۃ�;�u�-  SSSSS�8�2=  �����   �M;�vދE�H�E�3��}�-������<0u��+ȍE�P�uQW�D  ��;�t��X�E�H9E������|-;E}(:�t
�G��u��_��u�E�j�u���u��������u�E�jP�u���u�u�������M�_^3�[�j�����U��E��et_��EtZ��fu�u �u�u�u�u�&�����]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u������u �u�u�u�u�u�|�����]�U��j �u�u�u�u�u�u�^�����]�VW3���h��6�  ����(Y�r�_^�Vh   h   3�V�LF  ����tVVVVV�:  ��^�U����Ȗ�]�����]��E��u��M��m��]����]�����z3�@��3���h�� ���thЖP����tj ���������������̀zuf��\���������?�f�?f��^���٭^�������剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�������剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp���������۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-����p��� ƅp���
��
�t���������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�"D  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   �� ��   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z��,������������������   s��<���$������������������   v��4��jh0��  j�D  Y�e� �u�N��t/�������E��t9u,�H�JP�[���Y�v�R���Y�f �E������
   �  Ë���j�  Y����̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t����U��$X�����(  �`�3ŉ��  ���Vtj
��   Y�B  ��tj�B  Y�����   ���   ���   ���   �]|�ux�}tf���   f���   f�]pf�Elf�ehf�md����   ���  ���  ���   �E�  ���   �@�jP���   �E�j P�h����E����EЍE�j �E�  @�u��E��(��E�P�$�j�
  �QS�\$VW3�3�;���tG��r���w  Uj�BF  ��Y�1  j�1F  ��Yu�=���  ���   �?  h��  S���U�/<  ����tVVVVV��3  ��h  ���Vj ��� �4���u&hМh�  V��;  ����t3�PPPPP�3  ��V�F;  @��<Yv8V�9;  ��;�j���h̜+�QP��D  ����t3�VVVVV�v3  ���3�hȜSU�.D  ����tVVVVV�R3  ���4���SU�D  ����tVVVVV�03  ��h  h��U�+B  ���3j��0���;�t%���t j �D$P�4����6�:  YP�6U�,�]_^[Y�j��D  ��Ytj�D  ��Yu�=��uh�   �4���h�   �*���YY�U��QQSV3��E�F3�P�u��]���  �}�Y~���BWS� ��p<�f9^�F�|0v#Wh��`�����YYt�FC��(;�r���e� �E�_^[��V�5���58��օ�t!������tP�5�����Ѕ�t���  �&h�� �����t#�J�����th�V����t
�t$�ЉD$�D$^�j ����Y�V�5���58��օ�t!������tP�5�����Ѕ�t���  �&h�� �����t#�������th,�V����t
�t$�ЉD$�D$^��<�� V�5���8�����u�5���k���Y��V�5���@���^á�����tP�5���A���Y�Ѓ���������tP�D������  jhP��  h�� ��E�u�F\��3�G�~��t/������t&h��u���Ӊ��  h,��u��Ӊ��  �~pƆ�   CƆK  C� ��FhP�H�j�B  Y�e� �E�Fl��u���Fl�vl�j.  Y�E������   �  �j�1  Y�VW���5���������Ћ���uNh  j�  ����YYt:V�5���5������Y�Ѕ�tj V�����YY� ��N���	V�����Y3�W�L�_��^�V��������uj�  Y��^�jhp���  �u����   �F$��tP����Y�F,��tP����Y�F4��tP����Y�F<��tP�q���Y�FD��tP�c���Y�FH��tP�U���Y�F\=��tP�D���Yj��  Y�e� �~h��tW�P���u�� �tW����Y�E������W   j�  Y�E�   �~l��t#W�t-  Y;=�t��0�t�? uW�+  Y�E������   V����Y�  � �uj�  YËuj�  YÃ=���tLW�|$��u&V�5���58��օ�t�5���5�����Ћ�^j �5���5���`���Y��W����_������t	j P�@��Wh�� �����u	�����3�_�V�5�h\�W��hP�W�����hD�W�����h<�W����փ=�� �5@����t�=�� t�=�� t��u$�8�����D�������5������<���������   �5��P�օ���   �u  �5��������5�����������5�����������5����������������g  ��teh���5������Y�Ѓ�����tHh  j�  ����YYt4V�5���5�������Y�Ѕ�tj V�����YY� ��N��3�@��l���3�^_ËD$���������t$������5������h�   �Ѓ��hx�� ���thh�P����t�t$����t$�����Y�t$�T��j��  Y�j�  Y�V������t�Ѓ�;t$r�^�V�t$3����u���t�у�;t$r�^ËL$V3�;�u�  VVVVV�    �,  ��jX^á��;�tډ3�^ËD$V3�;�u��  VVVVV�    �s,  ��jX^�95��tۋ���3�^Ã=�� th���>  ��Yt�t$���Y�S���hD�h,��6�����YYuTVWh������� ��ƿ(�;�Ys���t�Ѓ�;�r�=� _^th��=  ��Ytj jj ��3��jh���  j�  Y3��}�3�C9�t~���E��9}u[�5�������E��5�����YY���u�9}�t&���u�;u�r�> t��>����;�t�W����Y����hT��H��2���Yh\��X��"���Y�E������   �} u(��j�  Y�u�����3�C�} tj�   Y��s  �j j�t$�������jj j �������V�������V�Q  V�=  V�)  V�&���V�|=  V�6  V����V�Y=  hS��K�����$���^�VW3��t$�]�������Yu'9�vV�X����  ;�v��������uɋ�_^�VW3�j �t$�t$��=  ������u'9�vV�X����  ;�v��������u���_^�VW3��t$�t$��>  ����YYu-9D$t'9�vV�X����  ;�v��������u���_^�jTh����	  3��}��E�P�d��E�����j@j ^V�@���YY;��  ���5p��   �0�@ ���@
�x�@$ �@%
�@&
�x8�@4 ��@����   ;�r�f9}��
  �E�;���   �8�X�;�E�   ;�|���E�   �[j@j ����YY��tV�M������p ��   �*�@ ���@
�` �`$��@%
�@&
�`8 �@4 ��@��;�r��E�9=p|���=p�e� ��~m�E����tV���tQ��tK�uQ�`���t<�u���������4���E� ���Fh�  �FP�/;  YY����   �F�E�C�E�9}�|�3ۋ���5�����t���t�N��r�F���uj�X�
��H������P�0������tC��t?W�`���t4�>%�   ��u�N@�	��u�Nh�  �FP�:  YY��t7�F�
�N@�����C���g����5p�\�3��3�@Ëe��E����������  �VW���>��t1��   �� t
�GP�h����@   ;�r��6�J����& Y�����|�_^�S3�9�VWu��"  �5��3�;�u����   <=tGV�m-  Y�t�:�u�jGW������;�YY�=��tˋ5��U�@V�<-  ��E�>=Yt/jU�Z���;�YY�tJVUP�-  ����tSSSSS�t%  �����8u��5������������   3�Y]_^[��5���h�����������U��Q�MS3�9EV���U�   t	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�#=  ��Yt��} t
�M��E�F�ۋU�Mt2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=����Pt#�><  ��Yt��M�E�F��M��E���<  ��YtF���UF�V�����t� B�U��M�����E��^[t�  ���U���S3�9�VWu�O   h  ��VS���4���;É5��t8�E�u�u��U��E�PSS�}������E���=���?sJ�M���sB�����;�r6P������;�Yt)�U��E�P�WV�}�������E���H����5��3�����_^[��QQ� �SUVW�=|�3�3�;�j]u-�׋�;�t� �   �"����xu	�ţ ��� �����   ;�u�׋�;�u3���   f9��t�f9u��f9u�=x�SSS+�S��@PVSS�D$4�׋�;�t2U�����;�Y�D$t#SSUP�t$$VSS�ׅ�u�t$�J���Y�\$�\$V�t����X;�t;�u��p���;��p���8t
@8u�@8u�+�@��U�Z�����;�YuV�l��D���UVW������V�l���_^][YY�VW������;ǋ�s���t�Ѓ�;�r�_^�VW������;ǋ�s���t�Ѓ�;�r�_^�U��QQV�E�3�P�u��u��z�����YtVVVVV�9!  ���E�P������YtVVVVV�!  ���}�^u�}�r3�@��jX��3�9D$j ��h   P������$�u3���}������lu$h�  ��  ��Yu�5$�����%$� ��3�@�U3�=luTS��W3�9-P~1V�5T��h �  U�v�����6U�5$��Ӄ�G;=P|�^�5TU�5$���_[�5$�����-$�]�U��QQV���������F  �V\�l�W�}��S99t��k����;�r�k��;�s99u���3���t
�X�ۉ]�u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   �`��=d����;�}$k��~\�d9 �=`��d�B߃�;�|�]�� =�  ��~du	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�øcsm�9D$u�t$P����YY�3�����h��d�5    �D$�l$�l$+�SVW�`�1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�������̃�S�\$ UV�s35`�W�����D$ �D$   �{t�N�38�����N�F�38������D$(�@f�  �k����L$0�T$�D$�L$ �S�t^�Dm �L��ɍ\���D$t��� 7  ���D$|DL�D$�����ù|$ t$����t�N�38�|����N�F�38�l����D$_^][����D$    �ƋL$(�9csm�u*�=h t!hh�,0  ����t�T$(jR�h���L$,�6  �D$,9hth`�W�Ջ��6  �D$,�L$�H����t�N�38������N�V�3:������K���P6  �{��P���h`�W�˺�����g6  ����U����`��e� �e� SW�N�@�;ǻ  ��t��t	�Уd��`V�E�P����u�3u����3�� �3����3��E�P����E�3E�3�;�u�O�@����u������5`��։5d�^_[��jhض�j���3��]3�;���;�u�c  �    WWWWW��  ������S�=lu8j��  Y�}�S�?  Y�E�;�t�s���	�u���u��E������%   9}�uSW�5$���������*����3��]�u�j�   Y�VW3��(��<�t�u��p��8h�  �0���a/  ��YYtF��$|�3�@_^Ã$�p� 3���S�h�V�p�W�>��t�~tW��W�Q����& Y������|ܾp�_���t	�~uP�Ӄ�����|�^[�U��E�4�p����]�jh������3�G�}�3�9$�u�����j�3���h�   �{���YY�u�4�p�9t���nj����Y��;�u��  �    3��Qj
�Y   Y�]�9u,h�  W�\.  YY��uW����Y�  �    �]���>�W�f���Y�E������	   �E������j
�*���Y�U��EV�4�p��> uP�$�����Yuj�{���Y�6���^]�h@  j �5$������TuËL$�%x� �%P �\3��X�`   @ËP�Tk����T$+P��   r	��;�r�3��U����M�AV�uW��+y�������i�  ��D  �M��I���M���  S�1��U�V��U��U����]ut��J��?vj?Z�K;KuB�� �   �s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J;։M�v��;�t^�M�q;qu;�� �   �s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���� �Ls%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   �x�����   �d�5��h @  ��H� �  SQ�֋d�x��   ���	P�x��@�d����    �x��@�HC�x��H�yC u	�`��x��x�ueSj �p�֡x��pj �5$����P�x�k��T+ȍL�Q�HQP�  �E���P;x�v�m�T�\�E�x��=d[_^�á`V�5PW3�;�u4��k�P�5TW�5$����;�u3��x�`�5P�Tk�5Th�A  j�5$���;ǉFt�jh    h   W���;ǉFu�vW�5$���뛃N��>�~�P�F����_^�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W�����u����   �� p  ;��U�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[��U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I��?�M�vj?Y�M��_;_uC�� �   �s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O��?�L1�vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���� �Ls�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N��?�]�K�vj?^�E���   �u���N��?vj?^�O;OuB�� �   �s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���� �Ls�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[��U����P�Mk�T������M���SI�� VW}�����M���������3���U��\����S�;#U�#��u
��;؉]r�;�u�T��S�;#U�#��u
��;ى]r�;�u[��{ u
���];�r�;�u1�T�	�{ u
��;ى]r�;�u�����؅ۉ]u3��	  S�@���Y�K��C�8�t�\�C�����U�t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��ɍy�>u;x�u�M�;du�%x� �M���B_^[�ËD$3�;͐�tA��-r�H��wjXË͔��D���jY;��#����������u���Ã���v�����u���Ã��V������L$Q�����Y��������0^ËD$�|���5|�������Yt�t$�Ѕ�Yt3�@�3��U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]Ã%H �O'  �H3��U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]�U��� S3�9]u ����SSSSS�    �  ������   �M;�V�ut!;�u�����SSSSS�    �  ������S����;ȉE�w�M�W�u�E��u�E�B   �u�u�P�u���'  ��;��t�M�x�E����E�PS�%  YY��_^[���t$j �t$�t$�t$�8������U���(  �������������5���=|�f���f���f�x�f�t�f�%p�f�-l������E ����E����E������������  ���������	 ����   �`��������d�������������j�H0  Yj �(�h���$��=�� uj�$0  Yh	 ����P�������������������U��W�}3�������ك��E���8t3�����_��-�  t"��t��tHt3�ø  ø  ø  ø  �SUVW�  ��U3��^WS�<����~�~�~3��~���� ���+Ɗ�CMu���  �   ��ANu�_^][�U��$d�����  �`�3ŉ��  SW�E�P�v������   ��   3����  @;�r�E���ƅ�   t+�]����;�w+�@P���  j R茽����C�C��u�j �v�E��vPW���  Pjj �Z4  3�S�v���  WPW���  PW�vS�?2  ��DS�v���  WPW���  Ph   �vS�2  ��$3��LE���t�L���  ���t�L ���  ��  �Ƅ   @;�r��M��  �E�����3�)E��U���  ЍZ ��w�L�р� ���w�L �р� ���  A;�rŋ��  _3�[�����Ŝ  ��jh�������������$��Gpt�l t�wh��uj ����Y�������j�g���Y�e� �wh�u�;5(�t6��tV�P���u�� �tV�~���Y�(��Gh�5(��u�V�H��E������   뎋u�j�.���Y�U���S3�S�M������������u���   �Đ8]�tE�M��ap��<���u���   ����ۃ��u�E��@���   ��8]�t�E��`p���[��U��� �`�3ŉE�S�]V�uW�h�����3�;��}u�������3��  �u�3�9�0���   �E��0=�   r����  �f  ����  �Z  ��P�Ȑ���H  �E�PW������)  h  �CVP趺��3�B��9U�{�s��   �}� ��   �u�����   �F����   h  �CVP�o����M��k�0�u���@��u��*�F��t(�>����E���,�D;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   ����j�C�C��4�Zf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�.����C�S��s3��{����95���b�������M�_^3�[諾����jh8������M���������}�������_h�u�����E;C�W  h   ����Y�؅��F  ��   �wh���# S�u�����YY�E�����   �u��vh�P���u�Fh= �tP�h���Y�^hS�=H����Fp��   �$���   j�����Y�e� �C����C����C���3��E��}f�LCf�E��@��3��E�=  }�L�� �@��3��E�=   }��  ��(�@���5(��P���u�(�= �tP诸��Y�(�S���E������   �0j�q���Y��%���u �� �tS�y���Y�����    ��e� �E�����Ã=� uj��V���Y��   3��SUV�t$���   3�;�Wto=��th���   ;�t^9(uZ���   ;�t9(uP�������   �0  YY���   ;�t9(uP�������   �#0  YY���   �ʷ�����   迷��YY���   ;�tD9(u@���   -�   P螷�����   ��   +�P苷�����   +�P�}������   �r��������   �=0�t9��   uP�.  �7�K���YYj�~P[��(�t�;�t9(uP�*���Y9o�t�G;�t9(uP����Y��Ku�V����Y_^][�SUV�t$W�=H�V�׋��   ��tP�׋��   ��tP�׋��   ��tP�׋��   ��tP��j�^P]�{�(�t	���tP�׃{� t
�C��tP�׃�Mu؋��   �   P��_^][�V�t$��tSUW�=P�V�׋��   ��tP�׋��   ��tP�׋��   ��tP�׋��   ��tP��j�^P]�{�(�t	���tP�׃{� t
�C��tP�׃�Mu؋��   �   P��_][��^Å�t7��t3V�0;�t(W�8�������YtV�R����> Yu��0�tV�x���Y��^�3��jhX������������$��Fpt"�~l t�����pl��uj �����Y��������j�#���Y�e� �Fl�=��i����E��E������   ��j� ���Y�u�ËD$����U��$X�����(  �`�3ŉ��  V���   ���   ���   �]|�ux�}tf���   f���   f�]pf�Elf�ehf�md����   ���  ���  ���   �E�  ���   �@�jP���   �E�j P�%����E��EЍE؃��E�  ��u��E����j ���(��E�P�$���u��uj�4%  Yh  ����P������  3�^�����Ũ  ��U���5���3�����Yt]��j��$  Y]�����U����u�M�迸���E����   ~�E�Pj�u�-  ������   �M�H���}� t�M��ap��Ã=�� u�D$����A���j �t$����YY�U���SV�u�M��E����]�   ;�sT�M胹�   ~�E�PjS�-  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�\-  ��YYt�Ej�E��]��E� Y������ *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�4'  ��$���o�����u�E���M�3��e���}� t�M��ap�^[�Ã=�� u�D$�H���w�� �j �t$�����YY�U���(�`�3ŉE�SV�uW�u�}�M�������E�P3�SSSSW�E�P�E�P�B7  �E�E�VP�,  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�g�����U���(�`�3ŉE�SV�uW�u�}�M��P����E�P3�SSSSW�E�P�E�P�6  �E�E�VP�M1  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�����������U��WV�u�M�}�����;�v;���  ��   r�=L tWV����;�^_u^_]�������   u������r*��$����Ǻ   ��r����$���$����$�h��$H#ъ��F�G�F���G������r���$���I #ъ��F���G������r���$���#ъ���������r���$���I ���������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�p�����$� �I �Ǻ   ��r��+��$�t�$�p�����F#шG��������r�����$�p�I �F#шG�F���G������r�����$�p��F#шG�F�G�F���G�������V�������$�p�I $,4<DLTg�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�p�������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�ËL$S3�;�VWt�|$;�w����j^�0SSSSS���������1�t$;�u��ًъ�BF:�tOu�;�u������j"Y�����3�_^[�U��MSV�u3�;�W�yu����j^�0SSSSS�M��������   9]v݋U;ӈ~���3�@9Ew�|���j"Y�����;��0�F~�:�t��G�j0Y�@J;��M;ӈ|�?5|�� 0H�89t�� �>1u�A��~W�f���@PWV�������3�_^[]�U��Q�U�BS��VW��% �  ��  #ωE�B��پ   �%�� �ۉu�t;�t�� <  �(��  �$3�;�u;�u�Ef�M�X��L��<  �]����������M��E���ΉH�u��P������Ɂ���  �։P�t�M�_^f�H[��U���0�`�3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���u�����f���6  �uЉC�E։�EԉC�E�P�uV������$��t3�PPPPP�������M�_�s^��3�[�W���������������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j�����Y�U��E�M%����#�������Vt1W�}3�;�tVV�@?  YY�����j_VVVVV�8��������_��u��P�ut	�?  ���?  YY3�^]�U������   �`�3ĉ�$�   �E�SV�u�HW�L$t+Ht$HtHtHtHHtHutj��   �hj�
j�j�j[Q�~WS�D  ����uG�E��t��t��t�d$P���L$P�F����\$@���L$PW�NQPS�D$P�D$$P�*D  ��h��  �t$�]F  �>YYt�=H� uV�-F  ��Yu�6��E  Y��$�   _^[3�������]ËD$�0��4��8��<�ËD$�l�V9Pt��k�t$��;�r�k�L$^;�s9Pt3���58������Y�j hx������3��}�}؋]��Lt��jY+�t"+�t+�td+�uD�L������}؅�u����a  �0��0��`�w\���`���������Z�Ã�t<��t+Ht�z����    3�PPPPP������뮾8��8���4��4��
�<��<��E�   P�����E�Y3��}���   9E�uj�����9E�tP����Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.�`��M܋d��`��9M�}�M�k��W\�D�E���腿����E������   ��u�wdS�U�Y��]�}؃}� tj �2���Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3��~����U��� SVW����3�9D��E��]��]�]���   h���̐��;��y  �5�h��W��;��c  P�_����$x�W�D���P�J����$d�W�H���P�5����L��E�P������YYtSSSSS�Q������}�u,hH�W��P� ���;�Y�T�th0�W��P����Y�P��P��M�;�ty9T�tqP�?����5T����2���;�YY��tV;�tR��;�t�M�Qj�M�QjP�ׅ�t�E�u3�E�P�*�����YtSSSSS�������}�r	�M    �D�M   �;�H�;E�t1P�Ľ��;�Yt&��;ÉE�t�L�;E�tP覽��;�Yt�u��ЉE��5D�莽��;�Yt�u�u�u�u����3�_^[�ËD$S3�;�VWt�|$;�w�o���j^�0SSSSS���������=�t$;�u��ً�8tBOu�;�t��
BF:�tOu�;�u��'���j"Y����3�_^[�U��SV�u3�9]Wu;�u9]u3�_^[]�;�t�};�w�����j^�0SSSSS����������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x�����n���j"Y���낋L$V3�;�|��~��u���^á�����^��7���VVVVV�    ����������^ËD$��t���8��  uP����Y������̋L$f�9MZt3�ËA<��8PE  u�3�f�x�����������̋D$�H<��ASV�q3҅�W�Dv�|$�H;�r	�X�;�r����(;�r�3�_^[���������������U��j�h��h��d�    P��SVW�`�1E�3�P�E�d�    �e��E�    h   �<�������tU�E-   Ph   �R�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]�jh������跼���@x��t�e� ���3�@Ëe��E������ʶ��������h�!����Y�X�ËD$�\�ËD$�`���t$�ؐ3�@� jhط�;���3��}��5`��"���Y��;�uS�E�P����Y;�tWWWWW��������}�t!hȥ� �;�th��P����;�u�)"V�W���Y�`��}��u�u�։E��/�E� � �E�3�=  �����Ëe�}�  �uj�L��e� �E������E�������jh���v����M3�;�v.j�X3���;E�@u�g����    WWWWW�������3���   �M��u;�u3�F3ۉ]���wi�=luK������u�E;Xw7j����Y�}��u�����Y�E��E������_   �]�;�t�uWS�D�����;�uaVj�5$�����;�uL9=��t3V����Y���r����E;��P����    �E���3��uj�J���Y�;�u�E;�t�    �������jh��X����]��u�u����Y��  �u��uS� ���Y�  �=l��  3��}�����  j����Y�}�S� ���Y�E�;���   ;5XwIVSP���������t�]��5V�����Y�E�;�t'�C�H;�r��PS�u��:���S������E�SP�������9}�uH;�u3�F�u������uVW�5$����E�;�t �C�H;�r��PS�u�����S�u��������E������.   �}� u1��uF������uVSj �5$��������u�]j�����YË}����   9=��t,V�Z���Y������������9}�ul����P����Y��_����   �����9}�th�    �q��uFVSj �5$��������uV9��t4V�����Y��t���v�V�����Y�����    3�������z����|�����u�l�������P�#����Y����U����u�M������E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap���jj �t$j ��������SVW�T$�D$�L$URPQQh,'d�5    �`�3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�=  �   �C�=  �d�    ��_^[ËL$�A   �   t3�D$�H3��Ϡ��U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j��<  3�3�3�3�3���U��SVWj j h�'Q�K[  _^[]�U�l$RQ�t$������]� jh8������e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E������U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�^�����t3�@�3�[�������L3��U��QV�uV��F  �E�F��Yu������ 	   �N ����-  �@t����� "   ��S3ۨt��^��   �N�����F�F����f��F�^�]�u,��D  �� ;�t�D  ��@;�u�u�OD  ��YuV� D  Yf�FW��   �F�>�H��N+�I;��N~WP�u��B  ���E��M�� �F����y�M���t���t�����������������@ tjSSQ�o;  #����t%�F�M��3�GW�EP�u�B  ���E�9}�t	�N �����E%�   _[^���A@t�y t$�Ix��������QP�z���YY���u	���U��V����M�E�M�����>�t�} �^]��G@SV����t4� u.�D$�-��L$������C�>�u������8*u�ϰ?�i����|$ �^[�U��$�����x  �`�3ŉ��  ��   S��  V3�W��  ��  �M��EЉ}ԉu��u�u��u��uĉu��u��"���9u�u-�|���VVVV�    V�������}� t�E��`p������  �E��@@��   P�CD  ���Yt6�u��5D  ���Yt(�u��'D  �u����4���D  ����YY3������@$�u����u���C  ���Yt6�u���C  ���Yt(�u���C  �u����4����C  ����YY3������@$��"���;������3Ʉ҉ủu؉u��U���  C�}� �]���  ��, <Xw����Х��3��3�3�����j��Y;��E��z  �$�!4�M���u��u��u��uĉu�u��X  �� t>��t-��tHHt���9  �M��0  �M��'  �M��  �M�   �  �M��	  ��*u ���}ԋ�;��}���  �M��]���  �E�k�
�ʍDЉE���  �u���  ��*u���}ԋ�;��}���  �M���  �E�k�
�ʍDЉE��  ��ItF��ht8��lt��w�x  �M�   �l  �;luC�M�   �]��W  �M��N  �M� �E  �<6u�{4uCC�M� �  �]��(  <3u�{2uCC�e�����]��  <d�  <i��  <o��  <u��  <x��  <X��  �u��E�P��P�u���  Y���E�Yt�MЍu�������C���]���  �MЍu�������  ��d�r  ��  ��S��   tZ��AtHHt@HHtHH�N  �� �E�   �U�M�@9u��]�   �]܉E���  �E�   �	  f�E�0uu�M�   �lf�E�0u�M�   �M����u������f�E��}ԋ��}���  ;�u�$��E܋E��E�   �  ��X�9  HHt]+��d���HH��  ��f�E��}�t'�G�Ph   �E�P�E�P��A  ����t�E�   ��G��E��E�   �E�E��P  ���;Ɖ}�t.�H;�t'f�E� � �M�t�+����E�   �  �u��  � ��E�P�'���Y��  ��p��  �t  ��e��  ��g�������itY��nt��o��  �E��E�   tI�M�   �@�7���}��?  ����  �E� t	f�E�f���Ẻ�E�   �  �M�@�E�
   �M�f���C  ��W���k  u��guG�E�   �>9E�~�E��}�   ~-�u���]  V�=������U�Y�E�t
�E܉u�����E�   3�����E��G��E��E�P�u����u��}�P�u��E�SP�5��襫��Y�Ћ}����   t9u�u�E�PS�5������Y��YY�}�gu;�u�E�PS�5���`���Y��YY�;-u�M�   C�]�S�r����E�   �M��!��s�p���HH��������Y  �E�'   �E��E�   ������E�Q�E�0�E��E�   ����f�� ��������� t��@�}�t�G���G�����@�G�t��3҉}���@t;�|;�s�؃� �ځM�   f�E� ��ڋ�u3ۃ}� }	�E�   ��e���   9E�~�E����u!Eč��  �E��M������t$�EؙRPSW�)0  ��0��9�]�����~M��N�̍��  +�Ff�E� �E؉u�tL��t�΀90tA�M܋M��0@�2If90t@@;�u�+E����;�u� ��E܋E��I�8 t@;�u�+E܉E؃}� ��   �E�@t%f� t�E�-��t�E�+��t�E� �E�   �]�+]�+]��E�u�uЍE�Sj �;������uċ}ЍE̍M��K����E�Yt�E�uWSj0�E��������}� �E�tQ��~M�u܉E���M�Pj���  P�E�FPF��=  ����u9E�t�u��E̍��  ������}� Yu���M����M�P�E������Y�}� |�E�tWSj �E��������}� t�u�規���e� Y�]�����E�t$�M��}Ԋ��)��������    3�PPPPP�$����}� t�E��`p��E̋��  _^3�[�������  ���-V,q,�,�,-9-1.�%D �U����`�3ŉE�SV3�9d�W��u8SS3�GWhL�h   S����t�=d������xu
�d�   9]~"�M�EI8t@;�u�����E+�H;E}@�E�d�����  ;���  ����  9] �]�u��@�E �5А3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w�.  ��;�t� ��  �P�Ԍ��;�Yt	� ��  ���E���]�9]��=  W�u��u�uj�u �օ���   �5�SSW�u��u�u�֋�;ˉM���   f�E t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w�Q-  ��;�tj���  ���P����;�Yt	� ��  �����3�;�tA�u�VW�u��u�u����t"9]SSuSS��u�u�u�VS�u �x��E�V����Y�u�������E�Y�Y  9]�]�]�u��@�E9] u��@�E �u�:  ���Y�E�u3��!  ;E ��   SS�MQ�uP�u ��:  ��;ÉE�tԋ5��SS�uP�u�u��;ÉE�u3��   ~=���w8��=   w�;,  ��;�t����  ���P�����;�Yt	� ��  �����3�;�t��u�SW袋�����u�W�u�u��u�u��;ÉE�u3��%�u�E��uPW�u �u��:  ���u������#u�W�����Y��u�u�u�u�u�u�����9]�t	�u�觋��Y�E�;�t9EtP蔋��Y�ƍe�_^[�M�3��2�����U����u�M��.����u(�M��u$�u �u�u�u�u�u�-����� �}� t�M��ap���U��QQ�`�3ŉE��h�SV3�;�W��u:�E�P3�FVhL�V����t�5h��4����xu
jX�h���h�����   ;���   ����   9]�]�u��@�E�5А3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w�X*  ��;�t� ��  �P����;�Yt	� ��  ���؅�ti�?Pj S�ĉ����WS�u�uj�u�օ�t�uPS�u���E�S�����E�Y�u3�9]u��@�E9]u��@�E�u��7  ���Yu3��G;EtSS�MQ�uP�u��7  ����;�t܉u�u�u�u�u�u��;��tV虉��Y�Ǎe�_^[�M�3��7�����U����u�M��3����u$�M��u �u�u�u�u�u�������}� t�M��ap���V�t$����  �v�/����v�'����v�����v�����v�����v�����6� ����v ������v$������v(�����v,������v0�؈���v4�Ј���v�Ȉ���v8������v<踈����@�v@譈���vD襈���vH蝈���vL蕈���vP荈���vT腈���vX�}����v\�u����v`�m����vd�e����vh�]����vl�U����vp�M����vt�E����vx�=����v|�5�����@���   �'������   �������   �������   �������   ��������   ��������   �������   �ڇ�����   �χ�����   �ć�����   蹇����,^�V�t$��t5�;��tP蛇��Y�F;��tP艇��Y�v;5��tV�w���Y^�V�t$��t~�F;��tP�Z���Y�F; �tP�H���Y�F;�tP�6���Y�F;�tP�$���Y�F;�tP����Y�F ;�tP� ���Y�v$;5�tV����Y^��U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^��U���S�u�M������]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�o   ��YYt�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�N����� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[��U����u�M��S����E�M����   �A% �  �}� t�M��ap���j �t$����YY�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  �������W�M�E�u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���58�N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r;�ur��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�4���+8�;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�58�N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��<�A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;0��<���   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�0��D��3�@�   �D��e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+<���M���Ɂ�   �ً@�]���@u�M�U�Y��
�� u�M�_[��U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  �������W�M�E�u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5P�N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r;�ur��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�L���+P�;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5P�N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��T�A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;H��T���   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�H��\��3�@�   �\��e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+T���M���Ɂ�   �ًX�]���@u�M�U�Y��
�� u�M�_[��U���|�`�3ŉE��ES3�V3��E��EF3�9]$W�E��}��]��u��]��]��]��]��]��]��]�u貶��SSSSS�    �J�����3��  �U�U��< t<	t<
t<uB��0�B���/  �$�O�Ȁ�1��wjYJ�݋M$�	���   �	:ujY������+tHHt����  ���jY�E� �  뢃e� jY뙊Ȁ�1���u�v��M$�	���   �	:uj�<+t(<-t$:�t�<C�<  <E~<c�0  <e�(  j�Jj�y����Ȁ�1���R����M$�	���   �	:�T���:��f����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�]���<+t�<-t��`����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*�<	�u��n���j�����J��M��Ȁ�1��wj	��������+t HHt���;���j�����M��jY�@���j�o����u���B:�t�,1<v�J�(�Ȁ�1��v�:�뽃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�[����B:�}��O����M��E�O�? t�E�P�u��E�P�'  �E�3Ƀ�9M�}��E�9M�uE9M�u+E=P  ��  =������  �����`;��E���  }�ؾ��E���`9Muf�M�9M���  �E��}���T�����u��q  k�Ƌ�f�; ��]�r��}�����M��u��]��]��S
�M�3��E��EԉE؉E܋¿�  3�#�#�% �  f����<
����  f�����  f������  f���?w3��EȉE���  f��uG�E����u�}� u�}� u	f!M���  3�f;�u!G�C���u9Ku9u�M̉MȉM��  !M��u��E�   �M��U�Ʌ҉U�~U�Lă��M��]��M��U���	�e� �ʋV��
;�r;�s�E�   �}� �^�tf��E��m��M��}� ��]�FF�E��M��}� ����  f��~;�E�   �u-�u؋M��e�������M����ʁ���  f���u؉M��f��M����  f��}B��������E�t�E��M܋]؋U��m�����ًM������N�]؉M�u�9u�tf�M�f�}� �w�Mԁ��� �� � u3�}��u*�e� �}��u�e� f�}���u	f�E� �G�f�E���E���E�f����u�sf�M�f�MċM؉MƋM���M�f�}��f����e� %   � ���e� �Ẽ}� �m����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W�M�_^3�[��x����&IzI�IJHJ�J�J�J�JYKNK�JU���t�`�3ŉE�S�]VW�u�}�f��U��ʸ �  #ȁ��  f�ɉ]��E���E���E���E���E���E���E���E���E���E���E���E�?�E�   �M�t�C-��C f�ҋu�}�u.��u*��u&f!;f;�����$ �C�C�C0�C 3�@��  f�����   �   �;�f� u��t��   @uh���Qf��t��   �u��u;h���;�u0��u,h���CjP�������3���tVVVVV�ƽ�����C�*h���CjP�������3���tVVVVV蚽�����C3��  �ʋ�i�M  �������Ck�M���������ىM�3�����ۃ�`;�f�U�u�}�f�E��M���  }���ۃ�`�M�;���  �E�T�˃������y  k�M�f�9 ��M�r��}ĥ��Eĥ�MƉE����y
�U�3��Ͼ�  3�#�#��E��E��E�E��� �  f;֍���  f;���  f=����  f=�?w3��E�E�E���  3�f;�u@�E����u9u�u9u�u	f�u���  f;�u$�U�@�B���u9ru92u�u�u�u��  �}�u��}��E�   �U��u�҅��u�~X�T��U��U����U��U��u��6����փe� �4;�r;�s�E�   �}� �}��w�tf��E��m��M��}� �GG�E��M��}� �}���  f��~;�E�   �u-�U��}�u��e������U�������  f���}�U��f��R��  f��}H�����҉U���E�t�E��U��}�u��m�������U�������M��}�U�uσ}� tf�M�f�}� �w�U����� �� � u3�}��u*�e� �}��u�e� f�}���u	f�E� �@�f�E���E���E�f=�sf�U�f�U��U�U�U���U�f�E��f��Ƀe� ��   ��� ���e� �M���k���3��M���f���?��  �H  �u��E��ы�3�#�#�� �  f;Ӎ<�E��E��E�E�����  f;���  f������  f���?w�E���  f;�uG�E����u9E�u9E�u	f�E���  f;�uG�E����u
9E�u9E�t��e� �E��E�   �U��u�҅��u�~R�u؍T��u��U��U��u��6��e� �֋p��;�r;�s�E�   �}� �X�tf� �E��m��M��}� �@@�E��M��}� ����  3�f;�~<�E�   �u.�U��]�u��e����ڋU����ց���  f;��]�U��f;�M����  f;�}B��������E�t�E��U��]�u��m�����ڋU������H�]�U�u�9E�tf�M�f�}� �w�U����� �� � u1�}��u(�}���E�uf�}����E�u	f�E� �G�f�E���E���E�f���rf�ىE�E�Ɂ�   ��� ���M�3��6f�E�f�E��E�E�E���E�f�}���f��Ɂ�   ��� ���M�E�E��E�U��M�f�
t2��M9E'f�" f�}� ��B����$ �B�B0�B ����jY9M~�M�u���j���?  f�E�[�E��}�M��e������E�����K�}�E�uڅ�}2�ށ��   ~(�E�}�M��m�������E������N���}�E�؋E@���Z�]��E���   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B�ҋ�tA�Eȍ0;։U�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K���K�K<5}�M��D�;9u	�0K;]�s�;]��E�sCf� �*؀��ˈX�D �E��M�_^3�[�Bp���À;0uK;�s�;ًE�s�f�  f�}� ��@���ʀ��� �P�0�@ �����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u�����   ^t   �3���t��   ��SVW�   t���t   ��t   ��t   ��   �   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#с�   ^[t��   t
;�u �  Ã�@�@�  Ã�SUVW��|$�\$3���tjZ��t����t����t���� t����t��   �ˋ��   #ǽ   �   t =   t=   t;�u��
����   #�t;�u��   ���   f�� t��   �t$(�L$$����#�#��;D$��   ���������D$�l$��|$�\$3���tjZ��t����t����t���� t����t��   �ˋ�#�t$=   t=   t;�u����   ���   #�t��   u��   ���   f�� t��   �T$�=L ��  �����\$�D$3���yj^f� t��f� t��f� t��f� t��f� t��   �Ƚ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #Ã�@t-�  t��@u��   ���   ���   ��#|$$��#��;�u���   �"���P�D$,�V  Y�\$(�D$(3҄�yjZ�   ��t��f� t��f� t��f� t���   ��t��   ��#�t"��    t�� @  t;�u��   ����#Ã�@t-�  t��@u��   ���   ���   �L$��3���� t   �_^][���U��E�MSVW3��x�E3ۉx�EC���xt�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�&  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP��  �EPSj �u���M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]�U��j �u�u�u�u�u�u�
�����]�U����ESV3ۋ���C��u�t�]tS�%  Y����  �t�Etj�  Y����w  ����   �E��   j��  �EY�   #�tT=   t7=   t;�ub��M��������{L�H��M�����{,����2��M�����z������M�����z�p���p���������   ���   �E��   3��t����W�}�����D��   ��E�PQQ�$��  �M��]��� �����������}�E�������T���]�����Au���3��E�����f�E�����;�}"+��]�t��u���m��]�t�M�   ��m�Hu���t�E����]��E������_tj�   Y�e���u��Et�E tj �x   Y���3���^��[�ËD$��t~���X���� "   ��L���� !   �3��Q��<$�$Y�Q�<$���$Y�U��Q��}��E�M#M��#E�����E�m�E���QQ�L$��t�-L��\$���t����-L��$������t
�-X��$���t	�������؛�� t���$�YY�jhX�蔍��3�9LtV�E@tH9d�t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%d� �e��U�E�������e��U�t������������������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ����������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� j
j �t$��  ��������������Q�L$+ȃ����Y��  Q�L$+ȃ����Y��  U��SVWUj j h�c�u�  ]_^[��]ËL$�A   �   t2�D$�H�3��_d��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h�cd�5    �`�3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y�cu�Q�R9Qu�   �SQ�p��SQ�p��L$�K�C�kUQPXY]Y[� ���U��QQ�EV�u�E��EWV�E��  ���;�Yu貚��� 	   �ǋ��J�u�M�Q�u�P���;ǉE�u����t	P褚��Y�ϋ�����������D0� ��E��U�_^��jhx��>�������u܉u��E���u�I����  �.���� 	   �Ƌ���   3�;�|;pr!�����8����� 	   WWWWW蝩�����ȋ��������������L1��u&�ޙ���8�ę��� 	   WWWWW�\�����������[P�s  Y�}���D0t�u�u�u�u�������E܉U���v���� 	   �~����8�M���M���E������   �E܋U�聉����u�  Y�U��$������  �`�3ŉ�  ��   V3�9�$  �E��u��u�u3���  ;�u'�����0����VVVVV�    苨��������  SW��  �����4�������ǊX$������u��]�t��u3��$  ����u&褘��3��0舘��VVVVV�    � ������0  �@ tjj j ��  �~�������  �N  ��Y�9  ��D��,  �5w���@l3�9H�E���P��4�M�������  3�9M�t����  ����]��E�3�9�$  �E��G  �E��E����=  ��u�3���
���E��ǃx8 t�P4��  ��	  �`8 j��  P�E��P�������Yt4�M�+��$  3�@;��V  j�E�SP��  �������  C�E��jS�E�P�  �������  3�PPj��  Qj�M�QP�u�C�E��x������v  j �E�PV��  P�E�� �4�,����I  �E��M��9u��E��>  �}� ��   j �E�Pj��  P�E�� ƅ  �4�,�����  �}���  �E��E��a<t<u�33�f��
��CC�E��u��M�<t<u9�u���  f;E�Y��  �E��}� tjXP�E���  f;E�Y��  �E��E���$  9E��H����  ���E��T4��D8�k  3ɋ��@��+  �ۋE��M���   9�$  �E��t  ��u��M��e� +M��E�;�$  s'�U��E��A��
u
�E�� @�E��@�E��}�   rы؍E�+�j �E�PS�E�P��4�,�����  �E�E�;���  �E�+E�;�$  r��  ���E���   9�$  ��  ��u��M��e� +M��E�;�$  s3�U��E��AAf��
u�E�f�  @@�E��E�f�@@�}��  rŋ؍E�+�j �E�PS�E�P��4�,����$  �E�E�;��  �E�+E�;�$  �p����  9�$  �2  �M��e� +M�j���  ^;�$  s,�U��u��f��
u
f�  �u�u�f�Ɓ}�R  r�3�VVh�  ��  Q���  +��+���P��PVh��  �x���;�tyj �E�P��+�P��5  P�E�� �4�,���t	u�;���	���E�;�G�E�+E�;�$  �E��6����0j �M�Q��$  �u��0�,���t�E��e� �E��	���E��}� u]�}� t'j^9u�u腓��� 	   荓���0�6�u�蔓��Y�+�u���D@t�E��8u3���N����    �V����  �����E�+E�_[��  3�^�[����  ��jh�������E���u�����  ������ 	   ����   3�;�|;pr!�����8�Ԓ��� 	   WWWWW�l������ɋ��������������L1��t�P�h  Y�}���D0t�u�u�u�?������E���q���� 	   �y����8�M���E������	   �E�胂����u�  Y��p�h   �bw����Y�L$�At�I�A   ��I�A�A�A   �A�a �ËD$���u����� 	   3��V3�;�|;pr�ґ��VVVVV� 	   �j�����3�^Ëȃ���������D��@^ø��á@��Vj^u�   �;�}�ƣ@jP��v����YY�8�ujV�5@��v����YY�8�ujX^�3ҹ����8���� ���� �|�j�^3ҹ��W�����������������t;�t��u�1�� B����|�_3�^��}  �=� t�R  �58��T��Y�V�t$���;�r"����w��+�����Q�7����N �  Y^Ã� V���^ËD$��}��P�����D$�H �  YËD$�� P���ËD$���;�r=��w�`���+�����P����YÃ� P���ËL$���D$}�`�����Q�ȃ��YÃ� P���ËD$V3�;�u����VVVVV�    膟�������^Ë@^á`���3�9t������U���SV�u3�;�W�}u;�v�E;�t�3���E;�t�������v�~���j^SSSSS�0���������R�u�M���W���E�9X��   f�Ef=� v6;�t;�vWSV�R�����/���� *   �$���8]�� t�M��ap�_^[��;�t.;�w(����j"^SSSSS�0蝞����8]�t��E��`p��u�����E;�t�    8]��0����E��`p��$����MQSWVj�MQS�]�p�x�;�t9]�b����M;�t�������z�H���;��k���;��c���WSV��Q�����S���j �t$�t$�t$�t$�������U����`�3ŉE�j�E�Ph  �u�E� �Ԑ��u����
�E�P����Y�M�3��V����U���4�`�3ŉE��E�M�E؋ES�EЋ V�E܋EW3�;E�M̉}��}��_  �5���M�QP�օ��Аt^�}�uX�E�P�u�օ�tK�}�uE�u܃���E�   u�u�跣����YF;�~[�����wS�D6=   w/������;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P��O��;�Yt	� ��  ���E���}�9}�t؍6PW�u��_P����V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u�x���t`�]��[9}ԋx�uWWWWV�u�W�u�Ӌ�;�t<Vj�r��;�YY�E�t+WWVPV�u�W�u��;�u�u��SP��Y�}���}��t�MЉ�u��?���Y�E��e�_^[�M�3���T����U����`�3ŉE��ESV3�9uW�E�N@  �0�p�p�F  ��X���}𥥥�����<�ыH�����Ή}���e� �������ˋ]���׍<;��0�P�Hr;�s�E�   3�9]�8t�r;�r��s3�C�ۉptA�H�H�U�3�;�r;�s3�F���Xt�@�M�H�e� �?�����<��P������Uމ�x�X��4;�U�r;�s�E�   �}� �0t�O3�;�r��s3�B�҉HtC�X�M�E�} �����3��&�H�����P�����������E���  �H�9ptջ �  �Xu0�0�x�E���  ������0�4?�H�����ʅˉp�Ht�f�M�f�H
�M�_^3�[�S����U��QQ�E�E�M�]��  ��������f�E��E���U�����U����Dz3��   3�f�E�uc�E�� u9MtU�]��������Au3�@�3���e�E   �t�M�eJ�Et�f�e��;�tf�M ��EQQQ�$�X������%Q���EQQ�$�C����U�����  �����  �E�]�U���VW�u�M��,R���E�u3�;�t�0;�u,�y���WWWWW�    �������}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP�����M������   ���B����t�G�ǀ�-u�M���+u�G�E���I  ���@  ��$�7  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   ���3��u���N��t�˃�0�f��t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �\�]��]ى]��G댨����u�u>��t	�}�   �w	��u,9u�v'�ۇ���E� "   t�M����E$�����ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^��U��3�9��P�u�u�uuh��P������]��Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ��L$S3�;�VW|[;psS������<���������@t5�8�t0�=��u+�tItIuSj��Sj��Sj�� ����3��趆��� 	   辆������_^[ËD$���u视���  茆��� 	   ����V3�;�|";ps�ȃ����������@u$�g����0�M���VVVVV� 	   ���������^Ë ^�jh���v���}����������4���E�   3�9^u6j
�z��Y�]�9^uh�  �FP荨��YY��u�]��F�E������0   9]�t������������D8P����E���u���3ۋ}j
�Py��YËD$�ȃ���������DP����U����`�3ŉE�V3�95��tN�=��u�Y  �����uf���pV�M�Qj�MQP����ug�=��u�����xuЉ5��VVj�E�Pj�EPV��P�x������t�V�U�RP�E�PQ����t�f�E�M�3�^�HM�������   ��U���SV�u3�;�t9]t8u�E;�tf�3�^[���u�M��M���E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P�|�����YYt}�E����   ��~%9M| 3�9]��R�uQVj	�p�А���E�u�M;��   r 8^t8]����   �e����M��ap��Y����ۃ��� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p�А���:����j �t$�t$�t$��������jhظ�is��3ۉ]�j� x��Y�]�j_�}�;=@}W�����8��9tD� �@�tP�  Y���t�E��|(�8���� P�h��8��4��F��Y�8��G��E������	   �E��%s���j�v��Y�SV�t$�F�Ȁ�3ۀ�u?f�t9�FW�>+���~,WPV����YP������;�u�F��y����F��N ���_�F�f �^��[�V�t$��u	V�3   Y^�V������Yt���^�f�F @tV�T���P�  YY���^�3�^�jh���&r��3��}�}�j�v��Y�}�3��u�;5@��   �8���98t^� �@�tVPV�i���YY3�B�U��8����H���t/9UuP�P���Y���t�E��9}u��tP�5���Y���u	E܉}��   F�3��u�8��4�V�h���YY��E������   �}�E�t�E��q���j�%u��Y�j����Y����������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��3�PPjPjh   @h������á����V�5�t���tP�֡����t���tP��^�SV�t$W3����;�u茀��WWWWW�    �$�������B�F�t7V����V����  V�]���P�  ����}�����F;�t
P�D��Y�~�~��_^[�jh ��p���M��3��u3�;���;�u�
����    WWWWW袏���������F@t�~�E��p���V����Y�}�V�/���Y�E��E������   �ՋuV�W���Y�jh@��o���E���u���� 	   ����   3�;�|;pr�y��� 	   SSSSS�������Ћ����<����������L��t�P����Y�]���Dt1�u����YP����u���E���]�9]�t����M���~��� 	   �M���E������	   �E��o����u�C���Y�V�t$WV�$������YtP����u	���   u��u�@Dtj�����j�������;�YYtV�����YP����u
�����3�V�E����������������Y�D0 tW�l~��Y����3�_^�jh`��!n���E���u�5~���  �~��� 	   ����   3�;�|;pr!�~���8��}��� 	   WWWWW芍�����ɋ��������������L1��t�P����Y�}���D0t�u�����Y�E���}��� 	   �M���E������	   �E��m����u�����Y�V�t$�F��t�t�v�2A���f����3�Y��F�F^����̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[��%ܐ������������h@��>��Y����̃=0� uK�(���t�$��Q<P�B�Ѓ��(�    �4���tV��蠇��V������4�    ^�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ĺ ں � �� � � &� 6� H� \� x� �� �� �� Ȼ ֻ � � �� � "� :� H� P� b� p� �� �� �� ̼ � �� � $� 2� @� Z� j� �� �� �� �� ֽ � �� � � 0� <� F� R� d� t� �� �� �� ľ Ծ � �� � � ,� <� N� ^� n� �� �� �� ��         0�        ]�� �(�m        �~�n            bad allocation  333333�?      �?               �H�����z>�@[ �� 0� �Q � �R P  [ pP ��  p �R `� p� �� �� �_ �� �_ �� PR �Z ` tool_KyamaSlide ...end Container Dump    - DA_MISSINGPLUG    - DA_CUSTOMDATATYPE     - DA_MARKER     - DA_ALIASLINK  - DA_CONTAINER  - DA_FILENAME (     - DA_STRING (  )    - DA_BYTEARRAY  - DA_LLONG  - DA_MATRIX     - DA_VECTOR     - DA_TIME   - DA_REAL   - DA_LONG   - DA_VOID  id:      - DA_NIL   Container Dump...             >@������.\source\KyamaSlide.cpp         ��������������   ����?-C��6?����MbP?      �?KyamaSlide_Tool.tif ...with enahncements by Keith Young - http://skinprops.com  KyamaSlide v1.3 - MultiSlide Tool by Anton Marchenko    ===========================================================     \�_ f:\maxon\cinema 4d r12\resource\_api\c4d_resource.cpp   #   M_EDITOR    ���� ��� <��� res     �������f:\maxon\cinema 4d r12\resource\_api\c4d_libs\lib_ngon.cpp  ���	�� г�� f:\maxon\cinema 4d r12\resource\_api\c4d_baseobject.cpp f:\maxon\cinema 4d r12\resource\_api\c4d_file.cpp   f:\maxon\cinema 4d r12\resource\_api\c4d_general.h  %s     f:\maxon\cinema 4d r12\resource\_api\c4d_basebitmap.cpp f:\maxon\cinema 4d r12\resource\_api\c4d_pmain.cpp  ���f:\maxon\cinema 4d r12\resource\_api\c4d_gv\ge_mtools.cpp   d��������0���Q�Q�@���    e+000      �~PA   ���GAIsProcessorFeaturePresent   KERNEL32                  �?5�h!���>@�������             ��      �@      �        runtime error   
  TLOSS error
   SING error
    DOMAIN error
  R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:    .mixcrt EncodePointer   KERNEL32.DLL    DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    CorExitProcess  mscoree.dll ����    	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ =    Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        ��������t�h�\�T�H�<����d�P�0��4�,��(�$� ������ ������������ܢآԢТ̢ȢĢ������������������������������t�l�`�H�<�(���ȡ����d�H�$��ܠ����������p�h�\�L�0�������l�P�,��ܞ�����GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL  InitializeCriticalSectionAndSpinCount   kernel32.dll    ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx                                                                                                                                                                                                                                                                                                ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun 1#QNAN  1#INF   1#IND   1#SNAN  _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   modf    fabs    floor   ceil    tan cos sin sqrt    atan2   atan    acos    asin    tanh    cosh    sinh    log10   log pow exp SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    CONOUT$     ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           `���              p�|���    �       ����    @   `��        ����    @   ��           ı��               ܱ�|���    4�       ����    @   ̱            X��           ,�@��|���    X�       ����    @   �            ���           ����    ��        ����    @   p�            ����           ȲԲ��    ��       ����    @   ��            ���           � ���    ��       ����    @   �            ��P�           `�l���    ��       ����    @   P�            ,���           ����    ,�        ����    @   ��            D��           �� ���    D�       ����    @   �            ��0�           @�H�    ��        ����    @   0�            ��x�           ����    ��        ����    @   x�            ����           дܴ��    ��       ����    @   ��            ��           �$�    �        ����    @   �            <�T�           d�l�    <�        ����    @   T�        �� ,' �c                     ����    ����    ����`�q�    ����    ����    ����    ��    ����    ����    ����     �    ����    ����    ����    ��    ����    ����    ����    3�    ����    ����    ����    �    ����    ����    ����    ������    ������    ����    ����    ;�    ����    ����    ��������    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����        ����    ����    ����    �
    ����    ����    ����    $    ����    ����    ����        ����    ����    �����!�!    ����    ����    �����!�!    ����    ����    �����"�"    ����    ����    ����    �#    ����    ����    ����    Z%    ����    ����    ����(((    ����    ����    ����b)b    ����    ����    ����    Ef    ����    ����    ����    Cm    ����    ����    ����    �y    ����    ����    ����    �|    ����    ����    ����    ~        �}����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    ���         Ŀ  �                     ĺ ں � �� � � &� 6� H� \� x� �� �� �� Ȼ ֻ � � �� � "� :� H� P� b� p� �� �� �� ̼ � �� � $� 2� @� Z� j� �� �� �� �� ֽ � �� � � 0� <� F� R� d� t� �� �� �� ľ Ծ � �� � � ,� <� N� ^� n� �� �� �� ��     FGetCurrentThreadId  GetCommandLineA HeapFree  �GetVersionExA HeapAlloc �GetProcessHeap  qGetLastError  �GetProcAddress  GetModuleHandleA  nUnhandledExceptionFilter  JSetUnhandledExceptionFilter �WriteFile �GetStdHandle  }GetModuleFileNameA  eTlsGetValue cTlsAlloc  fTlsSetValue dTlsFree ,InterlockedIncrement  (SetLastError  (InterlockedDecrement  � ExitProcess VSleep $SetHandleCount  fGetFileType �GetStartupInfoA � DeleteCriticalSection � FreeEnvironmentStringsA UGetEnvironmentStrings � FreeEnvironmentStringsW �WideCharToMultiByte WGetEnvironmentStringsW  HeapDestroy HeapCreate  �VirtualFree �QueryPerformanceCounter �GetTickCount  CGetCurrentProcessId �GetSystemTimeAsFileTime HeapSize  QLeaveCriticalSection  � EnterCriticalSection  �VirtualAlloc  HeapReAlloc ^TerminateProcess  BGetCurrentProcess 9IsDebuggerPresent GetCPInfo � GetACP  �GetOEMCP  ?IsValidCodePage RLoadLibraryA  uMultiByteToWideChar tGetLocaleInfoA  #InitializeCriticalSection �RtlUnwind DLCMapStringA  ELCMapStringW  �GetStringTypeA  �GetStringTypeW  �RaiseException  SetFilePointer  "GetConsoleCP  3GetConsoleMode  7SetStdHandle  �WriteConsoleA 5GetConsoleOutputCP  �WriteConsoleW S CreateFileA 4 CloseHandle � FlushFileBuffers  KERNEL32.dll                    �ՐN    �          � � � б !�   KyamaSlide.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       `���    .?AVToolData@@  ��    .?AVBaseData@@  ��    .?AVDescriptionToolData@@   ��    .?AVMSlide@@    `�`�`�`�`�`���    .?AVGeSortAndSearch@@   ��    .?AVTranslationMapNewSearch@@   ��    .?AVTranslationMapSearchN@@ ��    .?AVTranslationMapSearch@@  `�`�`�`�`���    .?AVNeighbor@@  ��    .?AVDisjointNgonMesh@@  `�`�`�`�`�`�`�`�`�`�`�`�`�`�`�`���    .?AVGeToolNode2D@@  ��    .?AVGeToolDynArray@@    ��    .?AVGeToolDynArraySort@@    ��    .?AVGeToolList2D@@  `�u�  s�      sqrt    `���    .?AVtype_info@@             N�@���D����������       ���5�h!����?      �?      `�                      p�   D�	   �
   ��   T�   $�    �   Ԛ   ��   t�   <�   �   ܙ   ��   X�     �!   (�"   ��x   x�y   h�z   X��   T��   D���������S�    �����
                                                                   �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �             x   
                                                                                                                                                                                                                                                                                                                      	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                                                                                                                                                                                                                                                                                     abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                      ��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    T�����C                                                                                              (�            (�            (�            (�            (�                              ��        P�ثX�0�0�   0� �        �إP�R���|�x�t�p�l�h�`�X�P�D�8�0�$� �������� ���������خЮ�Ȯ����������������x�d�X�	         0�.   ��l�l�l�l�l�l�l�l�l���   .         ���5      @   �  �   ����                h�   d�   `�   X�   P�   H�!   @�   8�   0�   (�    �   �   �   �    �   �   ��   ��   �   �   ܯ   ԯ   ̯   į"   ��#   ��$   ��%   ��&   ���&         �D        � 0              �            @�    @�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �p     ����    PST                                                             PDT                                                             �P�����        ����                 �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
          �      ���������              �           ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l      ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �                 0  �              	  H   X V   �      <assembly xmlns="urn:schemas-microsoft-com:asm.v1" manifestVersion="1.0">
</assembly>PAPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDING   �   Z0�0�0�0�01131C1a1�1�1212W2_2�2�2�2�2�23,3q3�3'4g4!5g5�5�5�5�5N6�67�7"9K9�9�9�:;<�<�=�=�=�=�=>2>C>c>�>�>�>�>?"?8?M?c?�?�?�?�?      ,  0)0?0]0o0�0�0�01181J1�1�1�1�1�12%2z2�2�2�2�2�23V3k3�3�3�3�3�304F4\4q4�4�4�45"575M5c5�5�5�5�56)6>6\6n6�6�67/7D7Z7p7�7�7�7�7�7�78�8�8�8�8�89929G9e9w9�9�9�9:":@:R:�:�:�:�:�:;1;F;O;d;y;�;�;�;�;�;�;<%<C<Y<s<�<�<�<�<�</=E=Z=c=x=�=�=�=�=�=	>>4>I>r>�>�>�>�>�>�>�>?&?/?F?]?t?�?�?�?�?�? 0  |    00,0R0e0w0�0�0�0�0�011'1H1L1P1T1X1\1`1d1h1l1p1t1x1|1:2Z2�2�3�3�3 4*4b4w4�4�4�425@5�5�5�5�5"606J89�:�;<�<w>�>   @  T   [0�01z1�1�1*2D2h2�2�2�2�2�2T3j3�3�3�4�4�5�587@7�8�89�9:.:Z:�<S=c=m=�=>3? P  �   601 1C1Q1d1w1�12�23:3m3�3�34J4�4�4�4�4%7A7�7�7>8|8�89�9�9�9�9�9:*:a:�:�:�:�:;;#;E;�;�;�;�;�;�;<<'<9<L<b<t<�<�<�<�<�<�<�<= =3=F=�=�=�=�=�=>>Q>d>�>�>�>�>�>?D?d? `     0401�1�122@2k2�3�3�3�34a4h4�4�45:5I5t5}5�5�5�5�5�5�5�566(6F6e6w6�6�6�6�6�67"7/7G7Y7k7}7�7�7�7�7�78848F8X8a88�8�8�8�8�8$929?9W9i9{9�9�9�9�9�9�9:(:D:V:h:q:�:�:�:�:�:;;-;N;d;�;�;�;�;�;�;<</<8<V<t<�<�<�<�<�<�<==@=V=r=�=�=�=�=�=�=>>;>W>i>�>�>�>�>?1?�?�?�?�?�?�?   p  �   0 010:0M0�0�0�01%1�1�1�1�1�1-2O2d2�2�2�2�2�2�263H3�3�34q4�4�4�455u5�5656u6�6�657�7�7%8e8�89U9�9�9E:�:�:5;�;�;<e<�<=U=�=�=E>�>�>5?�?�? �  l   %0u0�01e1�1�152u2�23e3�34U4�45U5�5�5E6�657�7�7%8u8�89e9�9:U:�:�:U;�;�;5<�<�<=�=�=!>q>�>!?q?�? �  �   0q0�01,1T1t1�122y2�2�23y3�3�3484\4x4�4�4�4=5U5�5,6Q6�6�6�6747T7a7�7�7�7�78t8949:4:T:�:�:�:;D;t;�;�;�;$<�<�<==="=)=0=7=>=H=R=Y=`=g=n=u=|=�=�=�=�=�=�=�=>9>�>e? �  $   �3a=�=�=�=%>e>�>�>5?r?�?�?   �  t   0R0�0�01E1�1�1�12B2u2�2�2E3�3�34U4�4�4E5�5�7�7P:�:�:�:�:�:�;�;�;�;r<�<�<�<n=|=�=�=�=�=�>
?#?1?�?�?�?�?   �  �   �0�0�0�01$1T1o1�1�1�1�12$2T2�2�2�2�2343d3�3�3�34$4Q4t4�4�4�4545T5t5�5�5�5�5616D6d6�6�6�6.7N7c7�78a8�8�8X9z9�9:::]:�:�:;~;�;�;3<\<�<�<�<$=�=�=>�>�>�>c?�?�? �  �   .0N0c0�0L1w1�1�1Q2w2�2�2Q3�334\4�4�4535�5�5�576�6�6l7�7�7�7�7�7$8D8[8�8�8�8�819Q9t9�9�9�9�9':Q:�:�:�:�:;+;J;�;�;�;�;<1<Q<t<====?=a=�=�=�=�=>$>T>�>�>�>�>?!?1?U?�?�? �  �    0.0g0�0�0�041d1�1�1�1�1!2D2a2�2�2�23$3T3�3�3�34b4�4�4�4�4545a5�5�5�5�5646d6�6�6�67$7D7d7�7�7�7�7818@8d8�8$9Q9d9�9�9�9:1:Q:�:�:�:�:;1;T;�;�;�;<D<t<�<�<=J=�=�=�=>!>D>t>�>�>�>�>�>?Z?t?�?�?   �  �   0:0�0�0�0�1�112E2Z2}2�2�2�233V33�3�34$4h4�4 5d5t5�5�5�5)6S6g6�6�6�6�6747d7�7�7�7�7848�8�8�8�8!9A9d9�9�9�9�9D:�:�:�:�:;_;~;�;�;<<H<c<�<�<�<�<=,=F=v=�=�=�=�=>?>S>h>�>�>�>?1?K?k?�?�?     �   Z0m0�0�0�0�0$1o1�3T6m6�6�677M7�7�7x9|9�9�9�9�9:1:B:d:u:�:�:�:�:�:�:;!;2;T;t;�;�;�;�;�;< <D<d<|<�<�<�<�<�<�<==/=@=}=�=�=�=�=�=>4>T>�>�>�>�>�>?$?T?t?�?�?�?�?    040Q0d0�0�0�0�011!141T1t1�1�1�1�1242T2t2�2�2�2�23�3(4:4O4p4x4�45?5[5q5�5�5�5646T6t6�6�6�6�6747T7q7�7�7�7�7�7�788,8T8s8�8�8�8�8�8!919A9Q9a9q9�9�9�9�9�9�9�9$:D:d:�:�:�:�:;$;D;w;�;�;�;�;�;<-<G<Y<�<�<�<�<=$=D=[=o=~=�=�=�=�=�=>>#>D>h>�>�>�>�>�>�>?!?2?T?r?�?�?�?�?     �   00D0Q0a0t0�0�0�0�0141T1t1�1�1�1�1242T2t2�2�2�2�2343T3|3�3�3�3444T4t4�4�4�4�4545T5t5�5�5�5�5646T6t6�6�6�6�6717D7d7�7�7�7�7�788$8D8d8�8�8�8�8�89:9t9�9�9�:�:�:�:�:2;G;�;�;�;�;!<4<d<�<�<�<�<$=T=t=�=�=>$>T>t>�>�>�>�>?4?F?a?t?�?�?�?�?�? 0 �   040q0�0�0�0�0141T1q1�1�1�1�1�12$2D2d2�2�2�2�2313D3d3�3�3�3�34T4z4�4�4�45$5D5d5�5�5�5�56D6�6�6�6C7�7�7�78D8q8�8�8�8�89!949T9t9�9�9�9	::r:�:�:�:;$;D;�;�;�;�;�;<&<6<d<�<�<�<�<=0=D=T=t=�=�=�=
>=>K>^>s>�>�>�>�>�>?"?2?T?x?�?�?�?�?   @ �   %0S0i0w0�0�0�0�0#191G1V1�1�1�1�1$2M2{2�2�2�23/3T3t3�3�3�3�34$4D4a4t4�4�4�4545T5t5�5�5�5�56!646Q6d6�6�6�6�6�67%767H7a7t7�7�7�78$8A8d8�8�8�8�8949Q9t9�9�9�9d:�:;$;D;a;t;�;�;�;<$<T<�<�<�<�<=J>\>n>�>p?w?~?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   P �   �0�1�1"2U2�2�23U3�3�3�3%4e4�4�4?5�5�5626e6�6�6B7u7�7858e8�8�89E9�9�9%:e:�:�:;0;D;T;u;�;<E<�<�<=U=�=�=>A>i>s>�>�>�>�>?E?i?�?�?   ` t   0/0�0�0�01=1f1�1�1262X2�23!3D3a3�3�3�3Q;d;�;�;�;�;<D<c<v<�<�<�<=A=T=�=�=�=�=>D>�>�>�>�>?T?t?�?�?�?�? p �   040d0�0�0�0Q1d1�1�1�12�3�3�3 4�45�6�6�6747T7�7�7�7�7�7�78D8t8�8�8�8�89$9A9d9�9�9�9�9�:;j;o;�;�<�<�<c=v=�=�=1>;>�>??4?T?t?�?�?�?�?   � �   0010A0T0q0�0�0�0�01(1A1d1�1�1�1�1242T2t2�2�2�2313A3T3t3�3�3�3�3414O4t4�4�4�4555M5\5�5�5�5�5�566-6q6�6�67K7�78U8�8�8&9u9�9�9(:�:�:;E;�;�;<X<�<�<"=U=�=�=�=E>�>�>�>�>
?2?u?�? � t   0R0�0�051�1�1%2r2�2�223u3�34�4�45�5�56V6�6�6E7�7�7(8�8(9�9�9%:b:�:�:E;�;�;%<u<�<=U=�=�=F>�>�>5?q?�?�?�? � �   E0�0�01e1�12e2�23e3�3�3%4f4�4�4E5�5�56o6�6�67\7�78|89Q9q9�9�9:T:�:�:;$;D;d;�;�;�;�;<$<T<t<�<�<�<=D=d=�=�=�=>?>a>�>�>�>?A?a?�?�?�?�? � �   0!0A0a0�0�0�0�01!1A1a1�1�1�1�1�1�1'2.2J2b2�2�2�2�2�2�2�2�2�23$3U3�3�3G4X4*8�8�8:P:�:�:�:;%;8;_;�;�;S<X<^<b<h<l<r<v<|<�<�<�<�<�<�<�<�<�<�<�<="=b=m==�=�=�=�= >&><>N>S>Y>_>�>�>�>�>�>�>�>>?D?_?�?�?�?   � �   0D0�0�001J1u1z1�1�1�1:2D2e2�2�23m33�3�3�3*4_4x44�4�4�4�4�4�45555555 5$5n5t5x5|5�5�5�56666 6A6k6�6�6�6�6�6�6�6�6�6
77777r7�78P8X8m8x8;�;�;   � �   	1�1`3�3�3�3�3�3�394�4H5�5{6|7�7�7�7�7�7�7�7�7�8�89�9�9�9�9:":F:O:V:_:�:�:�:�:;&;?;Q;v;�;�;<	<< <5<;<O<V<z<�<�<�<�<�<�<�<�<�<�<===!=-=;=A=M=S=`=j=p=}=�=�=�=�=�=�= >&>P>V>r>�>�>?=?G??�?�?�?�?�?�? � P  00"00070=0S0X0`0f0m0s0z0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 1111 1+101=1K1Q1a1~1�1�1�1�1�1�1�1�12�2�2�2�2�2�2333)303J3T3j3t3�3�3�3�3�3�3�34	4'4�4�4�4�4�45&525h5q5}5�5�5�5�56Y6a6�6�6�6�6-7]7o7�7�7�78)878F88�8�8�8�8�89�:�:�:�:�:�:H;N;a;k;�;�;�;�;�;,<><o<�<�<�<�<�<I=P=b=y==�=�=�=�=�=�=�=�=�=�=�=�=�=>�>�>�>�>�?�?�?   � �   �0�0�01`1}1�1�1�1�1�1�1�122E2�2�2�2�2�2�2�2�2"3)3B3T3Z3c3v3�3-4M4]4c4j4w4~4�4�4�4�4�4�6�6�677&7/7<7G7Y7l7w7}7�7�7�7�7�7�7�7�7�7�7�7�7�78888'848:8T8e8k8|8�8w<�<�<�<=[=.?9?A?\?w?�?�?�?�?     �   �0�083>3D3J3P3V3]3d3k3r3y3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�34	44%4,4�4 55~6�6�6�6�6�6�6767>7H7a7k7~7�7�788�8�8�8V9u9�9�9	::6:>:F:]:v:�:�:�:�:�:�:�:;;?;<*<t<�<�<B=�=�=�=
>5>I>�>�>�>??;?�?�?  �   �01�1�2�2�2�2�2�2�2�23C3a3h3l3p3t3x3|3�3�3�3�3�3�3�3F4Q4l4s4x4|4�4�4�4�45555555 5j5p5t5x5|5?8O:;C;H;M;R;];�;�;�;�;,<1<8<=<D<I<�<�<�<Z=q=w=�=�=�=�=�=�=�=�=>>>>,>:>�>�>�>     �   ?0F0L011-1K1_1e1�1222$2/2<2L2~2�2�2�2�2�2�23]3r3�3�3�34R4�4�4�4L5R5v5�5�5�5�5&6�6�6�7�7�8�9�9�:r;�;�;�;'<:<R<�>�? 0 p   �0�01�2!4%4)4-4145494=4C4P4_4o4{4�4�4�4�4�4�5>6a6�6�748>8V8]8g8o8|8�8�8L9�9�;�;�;<<(<:<L<^<p<�>z?�?   @ T   501�1�1X2^2n23%3�3�4�4w5Y6�6�6�7�7�7P8g8�8"9�;	<?"?&?*?.?2?6?:?>?B?F?J?U? P     +0C0R0~0�01�:i>�?�?�?   ` �   00�0�1�1�1�1�1�1.2�3�3�3q4�4�4�45595w5�5^6�6w7�7l8�8�8:�:d;�;�;�;�;t<�<�<O=�=�=�=�=>!>,>:>H>O>^>j>w>�>�>�>�>�>�>+?5?>?a?�?�?�? p �   �01T1q1�1�1�1�2�2M38.8z8�8�8�89&9`9|9�9�9::&:4:<:I:f:p:y:�:�:�:�:�:�:x;�;</<;<b<o<t<�<Q=t==�=�=�>�>�>�>�>�>b?�?   � 0   
020i0s0�011.1V1�1�1 313B3J3T3f3p3�3   � �   $1014181<1@1L1P1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1h4l4�4�4�4�4�4�45 5$5(5,5D6H6�6�6�6�6�6�6�6�6�6�6�6�=�=   � �   �3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5 �   T1X1l1p1t1|1�1�1�1�1�1�1�1�1�1�1222(2,2024282@2X2h2l2|2�2�2�2�2�2�2�2�2�2�2�2 3333 383H3L3\3`3d3l3�3�3�3�3�3�3�3�3�3�3�3�3 44(4,4<4@4H4`4p4t4�4�4�4�4�4�4�4�4�4�4�45555$5<5L5P5`5d5l5�5�5�5�56(6H6h6�6�6�6�6�6�6707P7p7�7�7�7�7�7�7�7808L8P8l8p8�8�8�8�89989X9x9 � |   00040X0p0t0x0|0�0�0�0�0�0�011 1$1(1,1D1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�12 282<2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�23333$3,343<3D3L3T3\3d3l3t3|3�3�3�3(; <�<�<�<�<�<�<�<�< ===== =$=(=,=0=4=8=<=@=D=H=L=P=T=X=\=`=d=h=l=p=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>>>> >d>l>t>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>????$?,?4?<?D?�?�?   �    �2�2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                