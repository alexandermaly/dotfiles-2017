MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       4�]�p�3�p�3�p�3��M�q�3�WN�h�3�W^��3г�n�s�3�p�2�&�3�W]�K�3�WI�q�3�WK�q�3�Richp�3�        PE  L ���O        � !  �  �      a     �                         �    
�                       � H   � (    P �                    ` 4                                  � @            �                            .text   ��     �                   `.rdata  8-   �  0   �             @  @.data    2                      @  �.rsrc   �    P     0             @  @.reloc  #   `  0   @             @  B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ��%V��H�QV�ҡ�%�T$�H�D$�IRj�PV�у���^� �����������́�   �L$�Q)  h���L$<�s)  h���L$�e)  �D$8P�L$Q��$�   R�N=  ��P�D$`P�`-  ��P�L$xQ�R-  ��P�L$ �-  �L$p��)  �L$T��)  ��$�   ��)  �$�)  �L$8�)  j j�j�j j ���T$L��R�])  hl� �'  ��4h���L$��(  h���L$<�(  �$P�L$<Q�T$xR�<  ��P�D$`P�,  ��P��$�   Q�,  ��P�L$ �e,  ��$�   �))  �L$T� )  �L$p�)  �L$8�)  �$�)  j j�j�j j ���T$L��R�(  hm� ��&  ��4�	  ��u�L$��(  3��Ĩ   á�%�H�A�$R�Ћ�%�Q�Jj j��D$hp�P�эT$R�^  ��%�H�A�T$R�Ѓ��L$�p(  �   �Ĩ   �����hl� �'  hm� ��&  ����������̋D$�� t ��t
-�  t3�ù�%�T  �����ø   �̡�%�D$�P�D$���   ���$P��� �������������̡�%�PH��p  j h�  Q�Ѓ�����̡�%�H@�T$�A,VR�������%�QQ���$�B,h�  ���Ћ�%�Q�B4jh�  ���и   ^� �����������̡�%SUVW�|$��H@�Q,W�ҋ\$�t$ ������   j ���h  � -�  to���  ��%���   �N�B��=)  u;��%���   �N�Pt�ҋء�%���   �Bt����;�u_�   �F^][� 3�_�F^]�   [� ��%���   �N�P��=2  uԡ�%���   �N�Bt�Ћ�%���   �؋Bt����;�u�_�   �F^][� ���F uK��%�Qj �ȋ��   h�  �Ѕ�u#�Qhm� �$  ����t_�   �F^][� �Rhl� ��VSW���Y  _^][� ��������̡�%SUVW�|$��H@�Q,W�ҋ\$��j �ˋ��Vg  � �����w'��%�P���   j h�  ����_��^�]��[� �L$$�T$ �D$QRPSW���{Y  _^][� ���̃���%�P�BlS�\$V�t$j Vh�  ���Ѕ��D$u^[��� W���z  �����|$u�G_^[��� ��%�Q�Blj Vh�  ���Ћ���u	_^[��� U����  ���t%���v  ���ky  ������  �u  ���D$ u]_^�   [��� ������$h�  �������\$3���~%�I �D� �D$������z
�L$ V��u  ��;�|ދ�%�Q���   jh�  ���Ћ�%�QH�t$$�D$���   h�  V�Ћ�%�QHj �苂p  h�  V�Ѓ�3ۅ����   ���%�Q\�J,P�D$$P3��у���t�   ��%�G�J\�T$ P�A,R�Ѓ���t���G��%�Q\�J,P�D$$P�у���t����%�G�J\�T$ P�A,R�Ѓ���t����;t$|
�L$S��t  ��;��[����L$ Q�\t  ��%���   �L$�P��j j��]_^3�[��� ���̡�%�P�Bl��V�t$ W�|$ j Vh�  ���Ѕ�u
_3�^��� ����w  ���D$u_�   ^��� ��%�Q�Blj Vh�  ���Ѕ��D$t�����}  ����tƋ�%�QH�t$(���   SUh�  V�Ћ�%�QH�؋��   h�  V�Ѓ��΋��������L$�t$0�Ԍ  j UVS�L$,���  ��t�=s  ���D$(u�L$輌  ][_�   ^��� ��    Qj W���  �L$ ���T$,R�D$P3�U�4t  ����   �D$��;D$,����   ���t0���N�Q�L$,�Cs  �V��L$(R�6s  ��L$(P�*s  �NQ�L$,�s  �V�������������F�����������������;Vt�F�������؃���;\$,~��t$0�L$,Q�L$�T$RU�ys  ���E����D$,P�L$Q�L$03�S�[s  ��tr��$    �t$��;t$,F�I ��%�D$    �Bl�L$0Q�L$$�T$R�PVQ�҃��|$0 t
���t$0����;t$,~��D$,P�L$Q�L$0S��r  ��u��T$(R�q  ��%���   �L$�B��j j�ЍL$��  ][_3�^��� �����������SUVW�|$������   �t$��t~�\$��tv��%���   �B����=�  u]��%�Q@�B,V�Ћ�����u
_�F^][� ��%�Q���   j h�  ���Ѕ�WS��Vu�{���_^][� ����_^][� _^]3�[� ��������������̡�%�H�A��$�T$VR�Ћ�%�Q�Jj j��D$$h��P�ы�%�B�P�L$Q�ҡ�%�H�Aj j��T$(hL�R�Ѓ�(�L$Q�L$�S  � j P�T$Rh� j	h'  �A  ��Phg� �6�  ���L$���hT  ��%�H�A�T$R�Ћ�%�Q�J�D$P�у���^��$����������V���P  �D$t	V�Y  ����^� ��Vh4�j4h�%j�,Z  ������t���LP  �����^�3�^���������������U��E��%� ]��U�졀%V��H�QV�ҡ�%�H�U�AVR�Ѓ���^]� U�졀%�P8�EPQ�JD�у�]� ���̡�%�H8�Q<�����U�졀%�H8�A@V�u�R�Ѓ��    ^]�������������̡�%�H8�������U�졀%�H8�AV�u�R�Ѓ��    ^]��������������U�졀%�P8�EP�EP�EPQ�J�у�]� ������������U�졀%�P8�EP�EPQ�J�у�]� ��%�P8�BQ�Ѓ����������������U�졀%�P8�EPQ�J �у�]� ����U�졀%�P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U�졀%�P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U�졀%�P8�EP�EPQ�J(�у�]� U�졀%�P8�EP�EP�EPQ�J,�у�]� ������������U�졀%�P8�EP�EP�EPQ�J�у�]� ������������U�졀%�P8�EP�EP�EP�EP�EPQ�J�у�]� ����U�졀%�P8�EP�EPQ�J0�у�]� U�졀%�P8�EP�EP�EPQ�J4�у�]� ������������U�졀%�P8�EPQ�J8�у�]� ����U�졀%�H��x  ]��������������U�졀%�H��|  ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H�A,]�����������������U�졀%�H�QV�uV�ҡ�%�H�Q8V�҃���^]�����̡�%�H�Q<�����U�졀%�H�I@]����������������̡�%�H�QD����̡�%�H�QH�����U�졀%�H�AL]�����������������U�졀%�H�IP]�����������������U�졀%�H��<  ]��������������U�졀%�H��,  ]��������������U�졀%�H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡�%�H���   �⡀%�H���  ��U�졀%�H�U�ER�UP�ER�UP���   Rh�.  �Ѓ�]����������������U�졀%�H�A]�����������������U�졀%�H��\  ]��������������U�졀%�H�AT]�����������������U�졀%�H�AX]�����������������U�졀%�H�A\]����������������̡�%�H�Q`����̡�%�H�Qd����̡�%�H�Qh�����U�졀%�H�Al]�����������������U�졀%�H�Ap]�����������������U�졀%�H�At]�����������������U�졀%�H��D  ]��������������U�졀%�H��  ]��������������U�졀%�H�Ix]�����������������U�졀%�H��@  ]��������������U��V�u���  ��%�H�U�A|VR�Ѓ���^]���������U�졀%�H���   ]��������������U�졀%�H��h  ]��������������U�졀%�H��d  ]��������������U�졀%�H���  ]�������������̡�%�H���   ��U�졀%�H��l  ]��������������U�졀%�H��   ]��������������U�졀%�H��  ]��������������U��V�u���B�  ��%�H���   V�҃���^]���������̡�%�H��`  ��U�졀%�H��  ]��������������U�졀%�H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U�졀%�H���  ]��������������U��U�E��%�H�E���   R���\$�E�$P�у�]�U�졀%�H���   ]��������������U�졀%�H���   ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H���   ]��������������U�졀%�H���   ]��������������U�졀%�H���   ]��������������U�졀%�H���   ]��������������U�졀%�H���   ]��������������U�졀%�H���   ]��������������U�졀%�P���E�P�E�P�E�PQ���   �у����#E���]����������������U�졀%�P���E�P�E�P�E�PQ���   �у����#E���]����������������U�졀%�P���E�P�E�P�E�PQ���   �у����#E���]����������������U�졀%�H��8  ]��������������U��V�u(V�u$�E�@��%�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@��%�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U�졀%�P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U�졀%�P0�EP�EP�EP�EPQ���   �у�]� ����̡�%�P0���   Q�Ѓ�������������U�졀%�P0�EP�EPQ���   �у�]� �������������U�졀%�P0�EP�EP�EP�EPQ���   �у�]� ����̡�%�P0���   Q�Ѓ������������̡�%�H0���   ��U�졀%�H0���   V�u�R�Ѓ��    ^]�����������U�졀%�H��H  ]��������������U�졀%�H��T  ]�������������̡�%�H��p  �⡀%�H���  ��U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H�U�E��X  ��VR�UPR�E�P�ыu�    �F    ��%���   �Qj PV�ҡ�%���   ��U�R�Ѓ� ��^��]��������U���$Vj hLGOg�M�躖  P�E�hicMCP�k������M����  ��%���   �JT�E�P�у���u(�u���Z�  ��%���   ��M�Q�҃���^��]á�%���   �AT�U�R�Ћu��P���Z�  ��%���   �
�E�P�у���^��]�������������U�졀%�H��  ]��������������U�졀%�H��\  ]��������������U�졀%�H�U��t  ��V�uVR�E�P�у����S  �M��  ��^��]�����U�졀%�H�U���  ��VWR�E�P�ы�%�u���B�HV�ы�%�B�HVW�ы�%�B�P�M�Q�҃�_��^��]����������������U�졀%�H�U���  ��VWR�E�P�ы�%�u���B�HV�ы�%�B�HVW�ы�%�B�P�M�Q�҃�_��^��]����������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H�U�E��VWj R�UP�ERP��t  �U�R�Ћ�%�Q�u���BV�Ћ�%�Q�BVW�Ћ�%�Q�J�E�P�у�(_��^��]��U�졀%�H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    ��%���   j P�BV�Ћ�%���   �
�E�P�у�$��^��]���U�졀%�H��8  ]��������������U���  ��3ŉE��M�EPQ������h   R� ����|	=�  |#���%�H��0  h\�hF  �҃��E� ��%�H��4  ������Rh���ЋM�3̓��l�  ��]�������U�졀%�H��  ��V�U�WR�Ћ�%�Q�u���BV�Ћ�%�Q�BVW�Ћ�%�Q�J�E�P�у�_��^��]����U�졀%�H��  ��V�U�WR�Ћ�%�Q�u���BV�Ћ�%�Q�BVW�Ћ�%�Q�J�E�P�у�_��^��]����U�졀%�H��p  ��$�҅�trh���M�虑  ��%�P�E�R4Ph���M��ҡ�%�P�E�R4Ph���M���j �E�P�M�hicMCQ������%���   ��M�Q�҃��M��t�  ��]�U�졀%�H��p  ��$V�҅�u��%�H�u�QV�҃���^��]�Wh!���M���  ��%�P�E�R4Ph!���M���j �E�P�M�hicMCQ������%���   �QHP�ҋu����%�H�QV�ҡ�%�H�QVW�ҡ�%���   ��U�R�Ѓ�$�M�譐  _��^��]������U�졀%�H��p  ��$V�҅�u��%�H�u�QV�҃���^��]�Wh����M���  ��%�P�E�R4Ph����M���j �E�P�M�hicMCQ������%���   �QHP�ҋu����%�H�QV�ҡ�%�H�QVW�ҡ�%���   ��U�R�Ѓ�$�M��ݏ  _��^��]������U�졀%�H��p  ��$�҅�u��]�Vh#���M��d�  ��%�P�E�R4Ph#���M���j �E�P�M�hicMCQ�������%���   �Q8P�ҋ�%���   ��U�R�Ѓ��M��E�  ��^��]���������������U�졀%�H��p  ��$�҅�u��]�Vhs���M��Ď  ��%�P�E�R4Phs���M���j �E�P�M�hicMCQ�W�����%���   �Q8P�ҋ�%���   ��U�R�Ѓ��M�襎  ��^��]���������������U�졀%�H���  ]��������������U�졀%�H��@  ]��������������U�졀%�H���  ]��������������U��V�u���t��%�QP��D  �Ѓ��    ^]������U�졀%�H��H  ]��������������U�졀%�H��L  ]��������������U�졀%�H��P  ]��������������U�졀%�H��T  ]��������������U�졀%�H��X  ]��������������U�졀%�H��\  ]�������������̡�%�H��d  ��U�졀%�H��h  ]��������������U�졀%�H��l  ]�������������̡�%�H���  ��U�졀%�H�U���  ��VR�E�P�ыu��P��蓌  �M�諌  ��^��]�����U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H���  ]��������������U�졀%�H��$  ]��������������U�졀%�H��(  ]��������������U�졀%�H��,  ]�������������̡�%�H��0  �⡀%�H��<  ��U�졀%�H���  ]�������������̡�%�H���  ��U�졀%�H���  ]������������������������������U�졀%�H��  ]�������������̡�%�H��P  �⡀%���   ���   ��Q��Y��������U�졀%�H�A�U��� R�Ћ�%�Q�Jj j��E�h��P�ыUR�E�P�M�Q�=   ��%�B�P�M�Q�ҡ�%�H�A�U�R�Ћ�%�Q�J�E�P�у�,��]��U�졀%�H�QV�uV�ҡ�%�H�U�AVR�Ћ�%�Q�B<�����Ћ�%�Q�M�RLj�j�QP���ҋ�^]���������h�%Ph�f 耋  ���������������U��h�%jh�f �\�  ����t
�@��t]�����]�������U��Vh�%jh�f �+�  ������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R�j  �E�NP�у�4�M���  ��^]ÍM�  ���^]��U��h�%jh�f 輊  ����t
�@��t]��3�]��������U��h�%jh�f 茊  ����t�x t�P]��3�]������U�졀%�P�EP�EP�EPQ�J�у�]� �����������̡�%V��H�QV�ҡ�%�H$�QDV�҃���^�����������U�졀%V��H�QV�ҡ�%�H$�QDV�ҡ�%�U�H$�AdRV�Ѓ���^]� ��U�졀%V��H�QV�ҡ�%�H$�QDV�ҡ�%�U�H$�ARV�Ѓ���^]� ��U�졀%V��H�QV�ҡ�%�H$�QDV�ҡ�%�H$�U�ALVR�Ѓ���^]� �̡�%V��H$�QHV�ҡ�%�H�QV�҃�^�������������U�졀%�P$�EPQ�JL�у�]� ����U�졀%�P$�R]�����������������U�졀%�P$�Rl]����������������̡�%�P$�Bp����̡�%�P$�BQ�Ѓ����������������U�졀%�P$��VWQ�J�E�P�ы�%�u���B�HV�ы�%�B�HVW�ы�%�B�P�M�Q�҃�_��^��]� ���U�졀%�P$�EPQ�J�у�]� ����U�졀%�P$��VWQ�J �E�P�ы�%�u���B�HV�ы�%�B$�HDV�ы�%�B$�HLVW�ы�%�B$�PH�M�Q�ҡ�%�H�A�U�R�Ѓ� _��^��]� ���U�졀%�P$��VWQ�J$�E�P�ы�%�u���B�HV�ы�%�B$�HDV�ы�%�B$�HLVW�ы�%�B$�PH�M�Q�ҡ�%�H�A�U�R�Ѓ� _��^��]� ���U���V�uV�E�P�l������e�����%�Q$�JH�E�P�ы�%�B�P�M�Q�҃���^��]� ����̡�%�P$�B(Q��Yá�%�P$�BhQ��Y�U�졀%�P$�EPQ�J,�у�]� ����U�졀%�P$�EPQ�J0�у�]� ����U�졀%�P$�EPQ�J4�у�]� ����U�졀%�P$�EPQ�J8�у�]� ����U�졀%�UV��H$�ALVR�Ѓ���^]� ��������������U�졀%�H�QV�uV�ҡ�%�H$�QDV�ҡ�%�H$�U�ALVR�Ћ�%�E�Q$�J@PV�у���^]�U�졀%�UV��H$�A@RV�Ѓ���^]� ��������������U�졀%�P$�EPQ�J<�у�]� ����U�졀%�P$�EPQ�J<�у������]� �������������U�졀%�P$�EP�EPQ�JP�у�]� U�졀%�P$�EPQ�JT�у�]� ���̡�%�H$�QX�����U�졀%�H$�A\]�����������������U�졀%�P$�EP�EP�EPQ�J`�у�]� �����������̡�%�H(�������U�졀%�H(�AV�u�R�Ѓ��    ^]��������������U�졀%�P(�R]����������������̡�%�P(�B�����U�졀%�P(�R]�����������������U�졀%�P(�R]�����������������U�졀%�P(�R ]�����������������U�졀%�P(�E�RjP�EP��]� ��U�졀%�P(�E�R$P�EP�EP��]� ��%�P(�B(����̡�%�P(�B,����̡�%�P(�B0�����U�졀%�P(�R4]�����������������U�졀%�P(�RX]�����������������U�졀%�P(�R\]�����������������U�졀%�P(�R`]�����������������U�졀%�P(�Rd]�����������������U�졀%�P(�Rh]�����������������U�졀%�P(�Rx]�����������������U�졀%�P(�Rl]�����������������U�졀%�P(�Rt]�����������������U�졀%�P(�Rp]�����������������U�졀%�P(�BpVW�}W���Ѕ�t:��%�Q(�Rp�GP���҅�t"��%�P(�Bp��W���Ѕ�t_�   ^]� _3�^]� ��U�졀%�P(�BtVW�}W���Ѕ�t:��%�Q(�Rt�GP���҅�t"��%�P(�Bt��W���Ѕ�t_�   ^]� _3�^]� ��U��VW�}W���0�����t8�GP���!�����t)�OQ��������t��$W��������t_�   ^]� _3�^]� ������������U��VW�}W���0�����t8�GP���!�����t)�O0Q��������t��HW��������t_�   ^]� _3�^]� ������������U�����%�E�    �E�    �P(�RhV�E�P���҅���   �E���uG��%�H�A�U�R�Ћ�%�Q�E�RP�M�Q�ҡ�%�H�A�U�R�Ѓ��   ^��]� ��%�Qh��h`  P���   �Ћ�%�����E��Q(u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P��-  ��3�^��]� �M��U�j ���Q�MR�����E�P�-  ���   ^��]� �������������U�졀%��V��H�A�U�R�Ѓ��M�Q��������^u��%�B�P�M�Q�҃�3���]� ��%�H$�E�I�U�RP�ы�%�B�P�M�Q�҃��   ��]� �U��Q��%�P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U�졀%�P(�R8]�����������������U�졀%�P(�R<]�����������������U�졀%�P(�R@]�����������������U�졀%�P(�RD]�����������������U�졀%�P(�RH]�����������������U�졀%�P(�E�R|P�EP��]� ����U�졀%�P(�RL]�����������������U�졀%�E�P(�BT���$��]� ���U�졀%�E�P(�BPQ�$��]� ����̡�%�H(�Q�����U�졀%�H(�AV�u�R�Ѓ��    ^]��������������U�졀%�P(���   ]��������������U�졀%�H(�A]����������������̡�%�H,�Q,����̡�%�P,�B4�����U�졀%�H,�A0V�u�R�Ѓ��    ^]�������������̡�%�P,�B8�����U�졀%�P,�R<��VW�E�P�ҋu����%�H�QV�ҡ�%�H$�QDV�ҡ�%�H$�QLVW�ҡ�%�H$�AH�U�R�Ћ�%�Q�J�E�P�у�_��^��]� �������U�졀%�P,�E�R@��VWP�E�P�ҋu����%�H�QV�ҡ�%�H�QVW�ҡ�%�H�A�U�R�Ѓ�_��^��]� ��̡�%�H,�j j �҃��������������U�졀%�P,�EP�EPQ�J�у�]� U�졀%�H,�AV�u�R�Ѓ��    ^]�������������̡�%�P,�B����̡�%�P,�B����̡�%�P,�B����̡�%�P,�B ����̡�%�P,�B$����̡�%�P,�B(�����U�졀%�P,�R]�����������������U�졀%�P,�R��VW�E�P�ҋu����%�H�QV�ҡ�%�H$�QDV�ҡ�%�H$�QLVW�ҡ�%�H$�AH�U�R�Ћ�%�Q�J�E�P�у�_��^��]� �������U�졀%�H��D  ]��������������U�졀%�H��H  ]��������������U�졀%�H��L  ]��������������U�졀%�H�I]�����������������U�졀%�H�A]�����������������U�졀%�H�I]�����������������U�졀%�H�A]�����������������U�졀%�H�I]�����������������U�졀%�H���  ]��������������U�졀%�H�A]�����������������U���V�u�E�P���������%�Q$�J�E�P�у���u-��%�B$�PH�M�Q�ҡ�%�H�A�U�R�Ѓ�3�^��]Ë�%�Q�J�E�jP�у���u=�U�R��������u-��%�H$�AH�U�R�Ћ�%�Q�J�E�P�у�3�^��]Ë�%�B�HjV�у���u��%�B�HV�у����I�����%�Q$�JH�E�P�ы�%�B�P�M�Q�҃��   ^��]�����������U�졀%�H�A ]�����������������U�졀%�H�I(]�����������������U�졀%�H��  ]��������������U�졀%�H��   ]��������������U�졀%�H��  ]��������������U�졀%�H��  ]��������������U�졀%�H�A$��V�U�WR�Ћ�%�Q�u���BV�Ћ�%�Q$�BDV�Ћ�%�Q$�BLVW�Ћ�%�Q$�JH�E�P�ы�%�B�P�M�Q�҃�_��^��]������U�졀%�H���  ��V�U�WR�Ћ�%�Q�u���BV�Ћ�%�Q$�BDV�Ћ�%�Q$�BLVW�Ћ�%�Q$�JH�E�P�ы�%�B�P�M�Q�҃�_��^��]���U�졀%�H���  ]��������������U���<��%��SVW�E�    t�E�P�   ��������/��%�Q�J�E�P�   �ы�%�B$�PD�M�Q�҃��}ࡀ%�H�u�QV�ҡ�%�H$�QDV�ҡ�%�H$�QLVW�҃���t)��%�H$�AH�U�R����Ћ�%�Q�J�E�P�у���t&��%�B$�PH�M�Q�ҡ�%�H�A�U�R�Ѓ�_��^[��]���U�졀%�H�U���  ��VWR�E�P�ы�%�u���B�HV�ы�%�B$�HDV�ы�%�B$�HLVW�ы�%�B$�PH�M�Q�ҡ�%�H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]���������̡�%�H���   ��U�졀%�H���   V�uV�҃��    ^]�������������U�졀%�P�]�⡀%�P�B����̡�%�P���   ��U�졀%�P�R`]�����������������U�졀%�P�Rd]�����������������U�졀%�P�Rh]�����������������U�졀%�P�Rl]�����������������U�졀%�P�Rp]�����������������U�졀%�P�Rt]�����������������U�졀%�P���   ]��������������U�졀%�P�Rx]�����������������U�졀%�P���   ]��������������U�졀%�P�R|]�����������������U�졀%�P���   ]��������������U�졀%�P���   ]��������������U�졀%�P���   ]��������������U�졀%�P���   ]��������������U�졀%�P���   ]��������������U�졀%�P���   ]��������������U�졀%�P���   ]��������������U�졀%�P���   ]��������������U�졀%�P���   ]��������������U�졀%�P���   ]��������������U�졀%�P�EPQ��  �у�]� �U�졀%�P���   ]��������������U�졀%�P���   ]��������������U�졀%�P���   ]��������������U��E��t ��%�R P�B$Q�Ѓ���t	�   ]� 3�]� U�졀%�P �E�RLQ�MPQ�҃�]� U��E��u]� ��%�R P�B(Q�Ѓ��   ]� ������U�졀%�P�R]�����������������U�졀%�P�R]�����������������U�졀%�P�R]�����������������U�졀%�P�R]�����������������U�졀%�P�R]�����������������U�졀%�P�R]�����������������U�졀%�P�E�R\P�EP��]� ����U�졀%�E�P�B ���$��]� ���U�졀%�E�P�B$Q�$��]� �����U�졀%�E�P�B(���$��]� ���U�졀%�P�R,]�����������������U�졀%�P�R0]�����������������U�졀%�P�R4]�����������������U�졀%�P�R8]�����������������U�졀%�P�R<]�����������������U�졀%�P�R@]�����������������U�졀%�P�RD]�����������������U�졀%�P�RH]�����������������U�졀%�P�RL]�����������������U�졀%�P�RP]�����������������U�졀%�P���   ]��������������U�졀%�P�RT]�����������������U�졀%�P�EPQ��  �у�]� �U�졀%�P���   ]��������������U�졀%�P���   ]��������������U�졀%�P�RX]����������������̡�%�P���   ��U�졀%�P���   ]��������������U�졀%�P���   ]��������������U�졀%�P���   ]��������������U�졀%�P���   ]�������������̡�%�P���   ��U�졀%�P���   ]�������������̡�%�P���   �ࡀ%�P���   �ࡀ%�P���   ��U�졀%�H���   ]��������������U�졀%�H��   ]��������������U�졀%�H�U�E��VWRP���  �U�R�Ћ�%�Q�u���BV�Ћ�%�Q�BVW�Ћ�%�Q�J�E�P�у�_��^��]������������U�졀%�H���  ]��������������U�졀%�P(�BPVW�}�Q�]���E�$�Ѕ�tM��%�G�Q(�]�E�BPQ���$�Ѕ�t,��%�G�Q(�]�E�BPQ���$�Ѕ�t_�   ^]� _3�^]� ����U�졀%�P(�BTVW�}����$���Ѕ�tE��%�G�Q(�BT�����$�Ѕ�t(��%�G�Q(�BT�����$�Ѕ�t_�   ^]� _3�^]� U��VW�}W��� �����t8�GP���������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U��VW�}W��� �����t8�GP��������t)�O0Q��������t��HW���������t_�   ^]� _3�^]� ������������U�졀%�} �P(�R8��P��]� ����U�졀%�P�BdS�]VW��j ���Ћ�%�Q�����   h����h�  V�Ћ�%�����Eu�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћ�%�Q(�BHV���Ѕ�t ��%�Q(�E�R VP���҅�t�   �3��EP�0  ��_��^[]� ����U���V�E���MP�K���P���#�����%�Q�J���E�P�у���^��]� ���U�졀%�P�E���   ��VWP�EP�E�P�ҋu����%�H�QV�ҡ�%�H�QVW�ҡ�%�H�A�U�R�Ѓ�_��^��]� ������������U��E��u��%�MP�EPQ�  ��]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3h��j;h�%j�  ����t
W���>����3����Fu_^]� �~ t3�9_��^]� ��%�H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   ��%�H<�Q��3Ʌ����^��������������̃y t�   ËA��uË�%�R<P��JP�у��������U����u��%�H�]� ��%�J<�URP�A�Ѓ�]� ���������������U�졈%��u��%�H�]Ë�%�J<�URP�A�Ѓ�]�U�졈%��$��Vu��%�H�1���%�J<�URP�A�Ѓ�����%�Q�J�E�SP�ы�%�B�P�M�QV�ҡ�%�H�A�U�R�Ћ�%�Q�Jj j��E�h�P�ы�%�B�@@�� j �M�Q�U�R�M��Ћ�%�Q�J���E�P���у���[t.��%�B�u�HV�ы�%�B�P�M�Q�҃���^��]á�%�P�E��RHjP�M��ҡ�%�P�E�M��RLj�j�PQ�M��ҡ�%�H�u�QV�ҡ�%�H�A�U�VR�Ћ�%�Q�J�E�P�у���^��]���������������U�졈%��$��SVu��%�H�1���%�J<�URP�A�Ѓ�����%�Q�J�E�P�ы�%�B�P�M�QV�ҡ�%�H�A�U�R�Ћ�%�Q�Jj j��E�h�P�ы�%�B�@@�� j �M�Q�U�R�M��Ћ�%�Q�J���E�P���у���t/��%�B�u�HV�ы�%�B�P�M�Q�҃���^[��]á�%�P�E��RHjP�M��ҡ�%�P�E�M��RLj�j�PQ�M��ҡ�%�H�A�U�R�Ћ�%�Q�Jj j��E�h�P�ы�%�B�@@��j �M�Q�U�R�M��Ћ�%�Q�J���E�P���у����3�����%�P�E��RHjP�M��ҡ�%�P�E�M��RLj�j�PQ�M��ҡ�%�H�u�QV�ҡ�%�H�A�U�VR�Ћ�%�Q�J�E�P�у���^[��]����������������U�졈%��$��SVu��%�H�1���%�J<�URP�A�Ѓ�����%�Q�J�E�P�ы�%�B�P�M�QV�ҡ�%�H�A�U�R�Ћ�%�Q�Jj j��E�h�P�ы�%�B�@@�� j �M�Q�U�R�M��Ћ�%�Q�J���E�P���у���t/��%�B�u�HV�ы�%�B�P�M�Q�҃���^[��]á�%�P�E��RHjP�M��ҡ�%�P�E�M��RLj�j�PQ�M��ҡ�%�H�A�U�R�Ћ�%�Q�Jj j��E�h�P�ы�%�B�@@��j �M�Q�U�R�M��Ћ�%�Q�J���E�P���у����3�����%�P�E��RHjP�M��ҡ�%�P�E�M��RLj�j�PQ�M��ҡ�%�H�A�U�R�Ћ�%�Q�Jj j��E�h�P�ы�%�B�@@��j �M�Q�U�R�M��Ћ�%�Q�J���E�P���у����������%�P�E��RHjP�M��ҡ�%�P�E�M��RLj�j�PQ�M��ҋu�E�P��������%�Q�J�E�P�у���^[��]�������U�졈%��$��SVu��%�H�1���%�J<�URP�A�Ѓ�����%�Q�J�E�P�ы�%�B�P�M�QV�ҡ�%�H�A�U�R�Ћ�%�Q�Jj j��E�h�P�ы�%�B�@@�� j �M�Q�U�R�M��Ћ�%�Q�J���E�P���у���t/��%�B�u�HV�ы�%�B�P�M�Q�҃���^[��]á�%�P�E��RHjP�M��ҡ�%�P�E�M��RLj�j�PQ�M��ҡ�%�H�A�U�R�Ћ�%�Q�Jj j��E�h�P�ы�%�B�@@��j �M�Q�U�R�M��Ћ�%�Q�J���E�P���у����3�����%�P�E��RHjP�M��ҡ�%�P�E�M��RLj�j�PQ�M��ҡ�%�H�A�U�R�Ћ�%�Q�Jj j��E�h�P�ы�%�B�@@��j �M�Q�U�R�M��Ћ�%�Q�J���E�P���у����������%�P�E��RHjP�M��ҡ�%�P�E�M��RLj�j�PQ�M���j h��M��R�����%�P�R@j �E�P�M�Q�M��҅���%�H�A�U�R���Ѓ���t/��%�Q�u�BV�Ћ�%�Q�J�E�P�у���^[��]Ë�%�M��B�PHjQ�M��ҡ�%�P�E�M��RLj�j�PQ�M��ҋu�E�P���˵����%�Q�J�E�P�у���^[��]���������������U�졀%�H<�A]����������������̡�%�H<�Q�����V��~ u>���t��%�Q<P�B�Ѓ��    W�~��t������W�d  ���F    _^��������U���V�E�P��������P��������M���i�����^��]��̃=�% uK��%��t��%�Q<P�B�Ѓ���%    ��%��tV��� ���V��  ����%    ^������������U���8��%�H�AS�U�V3�R�]��Ћ�%�Q�JSj��E�h�P�ы�%�B<�P�M�Q�ҋ�%�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��^  �M�Q�U�R�M��X^  ����   W�}�}���   ��%���   �U��ATR�Ћ�����tB��%�Q�J�E�P���у��U�Rj�E�P��������%�Q�ȋBxW�Ѕ��E�t�E� ��t��%�Q�J�E�P����у���t��%�B�P�M�Q����҃��}� u"�E�P�M�Q�M��]  ���;����E�_^[��]ËU��U�_�E�^[��]��������������U���DSV�u3�;�]�u_��%�H�A�U�R�Ћ�%�Q�JSj��E�h�P�ы�%�B<�P�M�Q�ҋ�%�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��\  �M�Q�U�R�M���\  ���p  W�}��I �E����   ��%���   �U��ATR�Ћ�������   ��%�Q�J�E�P���ы�%�B���   ���M�Qj�U�R���Ћ�%�Q�J���E�P�ы�%�B�P�M�QV�ҡ�%�H�A�U�R�Ћ�%�Q�Bx��W�M��Ѕ��Et�E ��t��%�Q�J�E�P����у���t��%�B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*��%���   P�BH�Ћ�%�Q���ȋBxW�Ѕ�t"�M�Q�U�R�M��r[  ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M���Z  �EP�M�Q�M�u��u�[  ����   �u���E���tA��t<��uZ��%���   �M�PHQ�ҋ�%�Q���ȋBxV�Ѕ�u-�   ^��]Ë�%���   �E�JTP��VP�[�������uӍUR�E�P�M��Z  ��u�3�^��]����������V��~ u>���t��%�Q<P�B�Ѓ��    W�~��t���j���W�$	  ���F    _^�������̋�� ��������������������̅�t��j�����̡�%�P��  �ࡀ%�P��(  ��U�졀%�P��   ��V�E�P�ҋuP�������M��������^��]� ��������̡�%�P��$  ��U�졀%�H��  ]��������������U�졀%�H���  ]�������������̡�%�H��  ��U�졀%�H���  ]��������������U�졀%�H��x  ]��������������U�졀%�H��|  ]��������������U���EV����t	V�  ����^]� �������������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������U���   V���_X  �����   �ESP�M��(�����%�Q�J�E�P�ы�%�B�Pj j��M�h��Q�҃��E�P�M������j j��M�Q�U�R��d���P������P�M�Q������P�U�R�������P�Y  ���M����!����M�������d��������M�������%�H�A�U�R�Ѓ��M��������[t	V�W  ����^��]� ���U��EVP����a  �����^]� �����Q�ZW  Y���������U��E�M�U�H4�M�P �U��M�@`l �@8`q �@<�q �@@�q �@D q �@H�q �@Lpq �@P0q �@l�q �@X r �@\@q �@`�q �@d�q �@T�q �@h�q �@pq �@tPq �P0�H(�@,    ]��������������U���   h�   ��`���j P贘  �M�U�Ej Q�MRPQ��`���R�����E �Uh�   ��`���Q�E��ERPj�%�����8��]��������������̋�`<����������̋�`����������̋�` ����������̋�`0����������̋�`@����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`����������̋�`����������̋�`,�����������U��V�u���t��%�QP��Ѓ��    ^]���������̡�%�H��@  hﾭ���Y����������U��E��t��%�QP��@  �Ѓ�]����������������U�졀%�H���  ]��������������U�졀%�H��  ]�������������̡�%�H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW���  ������u_^]Ã} tWj V�<�  ��_������F��%   ^]���U���%�ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW肛  ������u_^]�Wj V�ƕ  ��_������F��%   ^]�������������U���%�ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW��  ������u_^]�Wj V�F�  ��_������F��%   ^]�������������U���%�ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW肚  ������u_^]�Wj V�Ɣ  ��_������F��%   ^]�������������U���%�ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW��  ������u_^]�Wj V�F�  ��_������F��%   ^]�������������U��M��t-�=�% t�y���A�uP�g�  ��]á�%�P�Q�Ѓ�]��������U��M��t-�=�% t�y���A�uP�'�  ��]á�%�P�Q�Ѓ�]��������U�졀%�H�U�R�Ѓ�]���������U�졀%�H�U�R�Ѓ�]���������U���%�ɋEt#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   VW�xW辘  ������u_^]�Wj V��  ��_������F��%   ^]���������U���%�ɋEtL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËMQ������]�������U��E��w�   ��%��t�U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�ϗ  ������u_^]�Wj V��  ��_������F��%   ^]����������U��E��w�   ��%��t,�} �U�IR�URPt���   �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW�<�  ������u_^]�Wj V耑  ��_������F��%   ^]�������U�졀%�H�U�R�Ѓ�]���������U�졀%�H�U�R�Ѓ�]���������U�졀%�H�U�R�Ѓ�]���������U�졀%�H�U�R�Ѓ�]���������U�졀%�Hp�]�ࡀ%�Hp�h   �҃�������������U��V�u���t��%�QpP�B�Ѓ��    ^]���������U�졀%�Pp�EP�EPQ�J�у�]� U�졀%�Pp�EP�EPQ�J�у�]� U�졀%�Pp�EP�EPQ�J�у�]� U�졀%�Pp�EPQ�J�у�]� ����h�%PhD �`J  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d��������]� ���������U��h�%jhD �I  ����t
�@��t]��3�]��������Vh�%j\hD ���\I  ����t�@\��tV�Ѓ���^�����Vh�%j`hD ���,I  ����t�@`��tV�Ѓ�^�������U��Vh�%jdhD ����H  ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh�%jhhD ���H  ����t�@h��t
�MQV�Ѓ�^]� ������������Vh�%jlhD ���|H  ����t�@l��tV�Ѓ�^�������U��Vh�%h�   hD ���FH  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�%h�   hD ����G  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�%jphD ���G  ����t�@p��t�MQV�Ѓ�^]� ��%^]� ��U��Vh�%jxhD ���iG  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh�%j|hD ���)G  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh�%j|hD ����F  ����t�@|��t�MVQ�Ѓ������^]� �   ^]� ����������̋���������������h�%jhD �F  ����t	�@��t��3��������������U��V�u�> t+h�%jhD �SF  ����t�@��tV�Ѓ��    ^]�������U��VW�}����t0h�%jhD �F  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh�%jhD ����E  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh�%jhD ���E  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh�%j hD ���LE  ����t�@ ��tV�Ѓ�^�3�^���Vh�%j$hD ���E  ����t�@$��tV�Ѓ�^�3�^���U��Vh�%j(hD ����D  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh�%j,hD ���D  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh�%j(hD ���YD  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh�%j4hD ���D  ����t�@4��tV�Ѓ�^�3�^���U��Vh�%j8hD ����C  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh�%j<hD ���C  ����t�@<��t
�MQV�Ѓ�^]� ������������Vh�%jDhD ���LC  ����t�@D��tV�Ѓ�^�3�^���U��Vh�%jHhD ���C  ����t�M�PHQV�҃�^]� U��Vh�%jLhD ����B  ����u^]� �M�PLQV�҃�^]� �����������U��Vh�%jPhD ���B  ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh�%jThD ���lB  ����u^Ë@TV�Ѓ�^���������U��Vh�%jXhD ���9B  ����t�M�PXQV�҃�^]� U��Vh�%h�   hD ���B  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh�%h�   hD ���A  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh�%h�   hD ���fA  ����u^]� �M���   QV�҃�^]� �����U��Vh�%h�   hD ���&A  ����u^]� �M���   QV�҃�^]� �����U��Vh�%h�   hD ����@  ����u^]� �M���   QV�҃�^]� �����U��Vh�%h�   hD ���@  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh�%h�   hD �e@  ����u��%�H�u�QV�҃���^��]ËM���   WQ�U�R�Ћ�%�Q�u���BV�Ћ�%�Q�BVW�Ћ�%�Q�J�E�P�у�_��^��]��U��Vh�%h�   hD ����?  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�%h�   hD ���?  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�%h�   hD ���F?  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�%h�   hD ���?  ����t���   ��t�MQ����^]� 3�^]� �Vh�%h�   hD ����>  ����t���   ��t��^��3�^����������������U��Vh�%h�   hD ���>  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�%h�   hD ���6>  ����t���   ��t�MQ����^]� ��������U��Vh�%h�   hD ����=  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vh�%h�   hD ���=  ����t���   ��t��^��3�^����������������VW��3����$    �h�%jphD �_=  ����t�@p��t	VW�Ѓ����%�8 t����_��^�����U��SW��3�V��    h�%jphD �=  ����t�@p��t	WS�Ѓ����%�8 tsh�%jphD ��<  ����t�@p��t�MWQ�Ѓ������%h�%jphD �<  ����t�@p��t	WS�Ѓ����%V���7�����t���[����E��^t�8��~=h�%jphD �\<  ����t�@p��t	WS�Ѓ����%�8 u_�   []� _3�[]� ��������U��Vh�%j\hD ���	<  ����t3�@\��t,V��h�%jxhD ��;  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh�%j\hD ���;  ����t3�@\��t,V��h�%jdhD �;  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh�%j\hD ���F;  ����tG�@\��t@V�ЋEh�%jdhD �E��E�    �E�    �;  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh�%j\hD ����:  ����t\�@\��tUV��h�%jdhD �:  ����t�@d��t
�MQV�Ѓ�h�%jhhD �~:  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh�%j\hD ���9:  ������   �@\��t~V��h�%jdhD �:  ����t�@d��t
�MQV�Ѓ�h�%jhhD ��9  ����t�@h��t
�URV�Ѓ�h�%jhhD ��9  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh�%jthD ���9  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h�%j`hD �N9  ����t(�@`��t!�M�Q�Ѓ���^��]� �uh�%���_�����^��]� ������U���Vh�%h�   hD ����8  ����tR���   ��tH�MQ�U�R���ЋuP������h�%j`hD �8  ����t<�@`��t5�M�Q�Ѓ���^��]� �u�U�R���E�    �E�    �E�    ������^��]� �������������̡�%�H\�������U�졀%�H\�AV�u�R�Ѓ��    ^]�������������̡�%�P\�BQ�Ѓ���������������̡�%�P\�BQ�Ѓ����������������U�졀%�P\�EPQ�J�у�]� ����U�졀%�P\�EP�EPQ�J�у�]� U�졀%�P\�EPQ�J�у�]� ���̡�%�P\�BQ�Ѓ����������������U�졀%�P\�EPQ�J �у�]� ����U�졀%�P\�EP�EPQ�J$�у�]� U�졀%�P\�EP�EP�EPQ�J(�у�]� ������������U�졀%�P\�EPQ�J0�у�]� ����U�졀%�P\�EPQ�J@�у�]� ����U�졀%�P\�EPQ�JD�у�]� ����U�졀%�P\�EPQ�JH�у�]� ���̡�%�P\�B4Q�Ѓ����������������U�졀%�P\�EP�EPQ�J8�у�]� U�졀%�P\�EPQ�J<�у�]� ����U���SVW�}��j �ωu��������%�H\�QV�҃���S�������3���~?��I ��%�H\�U�R�U��EP�A(VR�ЋM��Q�������U�R��������;�|�_^[��]� �������������U���VW�}�E��P��������}� ��   ��%�Q\�BV�Ѓ��M�Q��������E���taS3ۅ�~L�I �UR�������E�P�������E;E�#����%�Q\P�BV�ЋE����;E��E~߃�;]�|�[_�   ^��]� _�   ^��]� �����������̡�%�PD�BQ�Ѓ���������������̡�%�PD�BQ�Ѓ���������������̡�%�PD�BQ�Ѓ����������������U�졀%�PX��Q�
�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ���������U�졀%�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U�졀%�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U�졀%�PX��`VWQ�J�E�P�ы��E���   ���_^��]� �������������U�졀%�PX�EPQ�J�у�]� ����U�졀%�PX�EPQ�J�у�]� ����U�졀%�PX�EPQ�J�у�]� ����U�졀%�PX�EPQ�J�у�]� ����U�졀%�PX�EPQ�J$�у�]� ����U�졀%�PX�EPQ�J �у�]� ����U�졀%�PD�EP�EPQ�J�у�]� U�졀%�HD�U�j R�Ѓ�]�������U�졀%�H@�AV�u�R�Ѓ��    ^]��������������U�졀%�HD�	]��U�졀%�H@�AV�u�R�Ѓ��    ^]��������������U�졀%�HD�U�j R�Ѓ�]�������U�졀%�H@�AV�u�R�Ѓ��    ^]��������������U�졀%�U�HD�Rh2  �Ѓ�]����U�졀%�H@�AV�u�R�Ѓ��    ^]��������������U�졀%�U�HD�RhO  �Ѓ�]����U�졀%�H@�AV�u�R�Ѓ��    ^]��������������U�졀%�U�HD�Rh'  �Ѓ�]����U�졀%�H@�AV�u�R�Ѓ��    ^]�������������̡�%�HD�j h�  �҃�����������U�졀%�H@�AV�u�R�Ѓ��    ^]�������������̡�%�HD�j h:  �҃�����������U�졀%�H@�AV�u�R�Ѓ��    ^]��������������U���3��E��E���%���   �R�E�Pj�����#E���]�̡�%�HD�j h�F �҃�����������U�졀%�H@�AV�u�R�Ѓ��    ^]�������������̡�%�HD�j h�_ �҃�����������U�졀%�H@�AV�u�R�Ѓ��    ^]��������������U��E����u��]� �E���%�E�    ���   �R�E�Pj������؋�]� ̡�%�PD�B$Q�Ѓ���������������̡�%�PD�B(Q�Ѓ���������������̡�%�PD�BQ�Ѓ���������������̡�%�PD�B(Q�Ѓ���������������̡�%�PD�BQ�Ѓ���������������̡�%�PD�B(Q�Ѓ���������������̡�%�PD�BQ�Ѓ���������������̡�%�PD�B(Q�Ѓ���������������̡�%�PD�BQ�Ѓ���������������̡�%�PD�B(Q�Ѓ���������������̡�%�PD�BQ�Ѓ���������������̡�%�PD�B(Q�Ѓ���������������̡�%�PD�BQ�Ѓ���������������̡�%�PD�B(Q�Ѓ���������������̡�%�PD�BQ�Ѓ���������������̡�%�PD�B(Q�Ѓ���������������̡�%�PD�BQ�Ѓ���������������̡�%�PD�B(Q�Ѓ���������������̡�%�PD�BQ�Ѓ����������������U�졀%�E�PH�B���$Q�Ѓ�]� ���������������U�졀%�PH�EPQ���   �у�]� �U�졀%�PH�EPQ���  �у�]� �U�졀%�PH�EPQ���  �у�]� �U�졀%�PH�EP�EPQ��  �у�]� �������������U�졀%�PH�EP�EPQ��  �у�]� ������������̡�%�PH���  Q�Ѓ�������������U�졀%�PH�EPQ���  �у�]� ̡�%�PH���   j Q�Ѓ�����������U�졀%�PH�EPj Q���   �у�]� ��������������̡�%�PH���   jQ�Ѓ�����������U�졀%�PH�EPjQ���   �у�]� ��������������̡�%�PH���   jQ�Ѓ����������U�졀%�PH�EPjQ���   �у�]� ���������������U�졀%�PH�EP�EPQ���   �у�]� �������������U�졀%�PH�EP�EPQ���   �у�]� ������������̡�%�PH���   Q�Ѓ�������������U�졀%�PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP���@���������t�E��%�QH���   PVW�у���_^]� �����U��EVW���MPQ�L���������t�M��%�BH���   QVW�҃���_^]� ̡�%�PH���   Q�Ѓ������������̡�%�PH���   Q�Ѓ�������������U�졀%�PH�EPQ���   �у�]� �U�졀%�PH�EPQ���   �у�]� �U�졀%�PH�EP�EPQ��8  �у�]� �������������U�졀%�PH�EP�EPQ��   �у�]� ������������̡�%�PH���  Q�Ѓ������������̡�%�PH���  Q�Ѓ������������̡�%�PH���  Q�Ѓ������������̡�%�PH��  Q�Ѓ������������̡�%�PH��  Q�Ѓ�������������U�졀%�PH�EP�EPQ��  �у�]� �������������U�졀%�PH�EP�EP�EPQ��   �у�]� ���������U�졀%�PH�EP�EP�EP�EPQ��|  �у�]� �����U�졀%�PH�EPQ��  �у�]� ̡�%�PH��T  Q�Ѓ�������������U�졀%�PH�EP�EPQ��  �у�]� �������������U�졀%�PH�EPQ��8  �у�]� �U�졀%�PH�EPQ��<  �у�]� �U�졀%�PH�EPQ��@  �у�]� �U�졀%�PH�EP�EP�EPQ��D  �у�]� ��������̡�%�PH��L  Q��Y��������������U�졀%�PH�EPQ��H  �у�]� ̡�%V��H@�Q,WV�ҋ�%�Q��j �ȋ��   h�  �Ћ�%�QH�����   h�  V�Ѓ���
��t_3�^Ë�_^�̡�%�P@�B,Q�Ћ�%�Q��j �ȋ��   h�  �������U�졀%�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U�졀%�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U�졀%�PH�EP�EP�EPQ��   �у�]� ��������̡�%�HH��  ��U�졀%�HH��  ]��������������U�졀%�E�PH��$  ���$Q�Ѓ�]� �����������̡�%�PH��(  Q�Ѓ�������������U�졀%�PH�EP�EPQ��,  �у�]� �������������U�졀%�E�PH�EP�E���$PQ��0  �у�]� ���̡�%�PH���  Q�Ѓ������������̡�%�PH��4  Q�Ѓ������������̋��     �������̡�%�PH���|  jP�у���������U�졀%�UV��HH��x  R��3Ƀ������^��]� ��̡�%�PH���|  j P�у��������̡�%�PH��P  Q�Ѓ������������̡�%�PH��T  Q�Ѓ������������̡�%�PH��X  Q�Ѓ�������������U�졀%�PH��Q��\  �E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����̡�%�PH��`  Q�Ѓ�������������U�졀%�PH�EPQ��d  �у�]� �U�졀%�E�PH��h  ���$Q�Ѓ�]� ������������U�졀%�E�PH��t  ���$Q�Ѓ�]� ������������U�졀%�E�PH��l  ���$Q�Ѓ�]� ������������U�졀%�PH�EPQ��p  �у�]� �U�졀%�PH�EP�EP�EP�EPQ���  �у�]� �����U�졀%�PH�EP�EP�EP�EP�EP�EPQ���  �у�]� �������������U�졀%�E�HH�U �ER�UP�E���$R�UP���   R�Ѓ�]������������U��U�E��%�HH�E���   R�U���$P�ERP�у�]����������������U���E�M�(��l  �M;�|�M;�~��]�����������U�졀%�PH�E���   Q�MPQ�҃�]� ������������̡�%�PH���   Q��Y�������������̡�%�PH���   Q�Ѓ������������̡�%�PH���   Q��Y��������������U�졀%�PH�EP�EPQ���   �у�]� �������������U�졀%�PH�EP�EP�EP�EP�EPQ���  �у�]� ̡�%�PH��t  Q��Y�������������̋�� 4��@    ��4���%�Pl�A�JP��Y��������U�졀%V��Hl�V�AR�ЋE����u
�   ^]� ��%�Ql�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uË�%�QlP�B�Ѓ�������U�졀%�Pl�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U��U�E��%�HH�ER�U���$P���  R�Ѓ�]����U�졀%�HH���  ]��������������U�졀%�HH���  ]��������������U��U0�E(��%�HH�E$R�U ���$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�,]������������U�졀%�HH���  ]��������������U�졀%�E�PH�EP���$Q���  �у�]� ��������U���SV���a����؅ۉ]���   �} ��   ��%�HH��p  j h�  V�҃����E�u
^��[��]� �MW3��}��p�������   �]��I �E�P�M�Q�MW�/�����tc�u�;u�[�I ������u�E�������L�;Ht-��%�Bl�S�@����QR�ЋD������t	�M�P������;u�~��}��M���}������;��r����]�_^��[��]� ^3�[��]� ����������U�����%SV�ًHH��p  j h�  S�]��ҋ�����u
^3�[��]� �E��u��%�HH���  �'��u��%�HH���  ���uš�%�HH���  S�ҋȃ��ɉEt�W������%�HH���   h�  S3��҃����  ���_�u����    ��%�Hl�U�B�IWP�ы�������   ��%�F�J\�UP�A,R�Ѓ���t�K�Q�M�������%�F�J\�UP�A,R�Ѓ���t�K�Q�M�����E��;Pt&�F��%�Q\�J,P�EP�у���t	�MS�l�����%�v�B\�M�P,VQ�҃���t�M�CP�C�����%�QH�E����   �E�h�  P�����у�;�����_^�   [��]� ������U�졀%�HH���   ]�������������̡�%�PH���   Q��Y��������������U�졀%�HH���  ]��������������U�졀%��P���   V�uW�}���$V�����E������At���E������z����؋�%�Q�B,���$V����_^]����������������U���0�%�U�V�u�U��]�W�P�}���   �E�PV�M�Q����� �@�@�E�����E��Au�����������z���������������z�����������Au������������z)���١�%�]��ɋ��]��]��P�RH�E�PV��_^��]���������Au������������������U�졀%�HH�]��U�졀%�H@�AV�u�R�Ѓ��    ^]�������������̡�%�HH�h�  �҃�������������U�졀%�H@�AV�u�R�Ѓ��    ^]��������������U�졀%�HH�Vh  �ҋ�������   �EPh�  ��������t]��%�QHj P���   V�ЋMQh(  �V�������t3��%�JH���   j PV�ҡ�%���   �B��j j���Ћ�^]á�%�H@�QV�҃�3�^]�������U�졀%�H@�AV�u�R�Ѓ��    ^]��������������U�졀%�HH�Vh�  �ҋ�����u^]á�%�HH�U�E��  RPV�у���u��%�B@�HV�у�3���^]�������U�졀%�H@�AV�u�R�Ѓ��    ^]��������������U�졀%�HH�I]�����������������U�졀%�H@�AV�u�R�Ѓ��    ^]��������������U�졀%�PH�EPQ���  �у�]� �U�졀%�PH�EPQ���  �у�]� ̡�%�PH���  Q�Ѓ�������������U�졀%�HH���  ]��������������U�졀%�E�HH�U0�E,R�U(P�E$R�U P�ER�U���\$�E�$P��P  R�Ѓ�,]������������̡�%�PH���  Q�Ѓ�������������U�졀%�PH�EP�EPQ���  �у�]� ������������̡�%�PH��  Q�Ѓ�������������U�졀%�PH�EP�EP�EPQ���  �у�]� ��������̡�%�PH���  Q�Ѓ������������̡�%�PH���  Q�Ѓ�������������U�졀%�PH�EPQ��  �у�]� �U�졀%�PH�EPQ��  �у�]� ̋������������������������������̡�%�HH���  ��U�졀%�HH���  ]��������������U�졀%�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ���������U�졀%�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ��������̡�%�PH��,  Q�Ѓ�������������U�졀%�PH�EPQ��X  �у�]� ̡�%�PH��\  Q�Ѓ�������������U�졀%�HH��0  ]��������������U�졀%��W���HH���   j h�  W�҃��} u�   _��]� Vh�  �������������   ��%�HH���   j VW�҃��M���  ��%�P�E�R0Ph�  �M����E��%�P�B,���$h�  �M��Ћ�%�Q@�J(j �E�PV�у��M���  ^�   _��]� ^3�_��]� �����U��S�]�; VW��u7��%�U�HH���   RW�Ѓ���u��%�QH���   jW�Ѓ���t�   �����   ��%�QH���   W�Ѓ��} u(��%�E�QH�M���  P�ESQ�MPQW�҃��B�u��t;��%�U�HH�ER�USP���  VRW�Ћ�%���   �B(�����Ћ���uŃ; u��%�QH���   W�Ѓ���t3���   ���Wu1��%�QH���   �Ћ�%�E�QH���   PW�у�_^[]� ��%�BH���   �у��} u0��%�M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� ��%�QH�h  �Ћ؃���u_^[]� ��%���   �u�Bx���Ћ�%���   P�B|���Ѕ�tU��%�E�QH�MP�Ej Q���  VPW�у���t��%���   �ȋBHS�Ћ�%���   �B(���Ћ���u�_^��[]� ��������������U��E��V��u��%�HH���  �'��u��%�HH���  ���u��%�HH���  V�҃���u3�^]� P�EP���>���^]� ���������U���D��%�HH���   S�]VWh�  S�ҋ�%�HH���   3�Wh�  S�u܉}��҃�;��E�}�}��}��p
  ��%���   �B����=�  ��%�  �QH���   Wh:  S�Ћ�%�QH�E����   h�  S�Ћ�%�QHW�����   h�  S�uԉ}��Ћ�%�QH�E苂  S�Ћ�%�QH�EЋ��  S�Ѓ�(���E��E�@��}   �M���M�MЅ�tMj�W�:  ���t@�@�Ẽ|� �4�~����%�������;�u/���C  ;E�~�E؋��pC  E���E�;Pu�E���E��E���;}�|��}� tv�u�j S�����������  ���������tV�������}�;�uK��%�H���  �4�hD���h�  V�҃����E��k  �M�PVP����P�$J  ����}ܡ�%�H���  �4�hD���h�  V�҃����E��   �M�3�;�t;�tVQP��Y  ���E�;�~-��%�QhD���h�  P���   �Ѓ�;ǉE���  ��%�E��QH��  j�PS�у�����  �u�;�tjS�����������  ��������E���}��%�BH���   Wh�  S�у�3�9}ԉE�}���  �}���}ȋMЅ��p  �U�j�R�8  ����\  �M̍@�|� ���]�~����%�������9E��  ���{A  �E�3�3�9C�E܉M���   ��I �����������t{�]��}������������ϋ9�<��}����҉��y�]��|��]������z�<��y�]��|��]������z�<��I�}��]������M��}ȃ��������M؃�;K�M��b������E��O  �+U�j��PR�M��#%  �M�v���E�3�+��U��E����	��$    ���E�;E���   �}� �U����E�t6�U�@�U�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�M��E�;]؍@�E��Ћ��P�Q�P�Q�P�Q�P�Q�@�A}c�UȋE�9�uX�ȋL�����������w4�$��� �U����4�"�M����t��U����t�
�M����t�M���;]�|��E�����;]؉M������U�;U��  �U�R�ѷ���E�P�ȷ���M�Q迷����_^3�[��]Ë�M�3�;G�Å���   �E�v�ЋW��R�ы��Q�P�Q�P�Q�P�Q�P�I�H�O��I�M�ы�P�Q�P�Q���ۉP�Q�P�Q�P�I�H��@�E�ЋU�Lv�ʋ��P�Q�P�Q�P�Q�P�Q�@�At8�G�U�@�ʋU�Lv	�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��w��U��@�ʋU���v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��w��U����@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�7����t?�G�U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�w�����O�E�����;EԉE��}�������U�R觵���E�P螵�����$  ���   �B����=  �  ��%�QH���   j h(  S�Ћ�%�QH�����   h(  S�ЋЃ�3��҉U�~#���ǅ�t�|� t�4N��tN���;�|�u��u܋�%�Q���  �4v�hD���hK  V�Ѓ����E���   �M��t��tVQP��S  ���u؋�%�Q���  �hD���hP  V�Ѓ����E�tP��t��tVWP�S  ���M����+�%�RH��PQ�E���   S�Ѓ���u�M�Q�\����U�R�S�����_^3�[��]á�%�HH���   j h�  S�҉E���%�HH���   j h(  S��3�3���3�9]؉E��}ĉ]��N  �U���    �څ��+  ���E�    ��   �U�<��v��   ����U��:��\:�Y�\:�Y�\:׉Y�Z�Y�R�Q�U��\�E��Y�\�T���Y�Z�Y�Z�Y�Z�Y�R�]��Q�U�����������;�|��}ă|� �w   �U��Eԍ8�I�ʋU�v���A�B�A�B�A�B�A�B�I�J�E���ЋE���v�Ћ��A�B�A�B�A�B�A�B�I�J�U���<ډ}ă�;]؉]�������M�3�3�;�~"�U����$    �d$ �t���   ��;�|�U�R�u������E�P�i�����_^�   [��]Ë�ܹ � � �� ��������U��E� �M+]� ���������������U��V��V�4���%�Hl�AR�Ѓ��Et	V�4�������^]� ���������̸   � ��������3�� �����������3�� �����������U��j P�EQRPV�~�����ǆ�   `� ǆ�   p� ǆ�   P� ]������������U�졀%�P�B<��   V�uW���Ѕ��}tj VW�Ӛ������u_^��]�h   ������j Q�H  �U �E�Mj R�UPQR������P�����Uh   ������QRWj�E�`� �E�p� �E�P� ��_����8_^��]���������������̋�`L����������̋�`D����������̋�`H����������̡�%�P�BVj j����Ћ�^���������U�졀%�P�E�RVj P���ҋ�^]� U�졀%�P�E�RVPj����ҋ�^]� ��%�P�B�����U�졀%�P���   Vj ��Mj V�Ћ�^]� �����������U�졀%�P�EPQ�J�у�]� ����U�졀%�P�EPQ�J�у������]� �������������U�졀%�P�E�RtP�ҋ�%���   P�BX�Ѓ�]� ���U�졀%�P�E�Rlh#  P�EP��]� ���������������U�졀%�P�E�RlhF  P�EP��]� ���������������U�졀%�P�E�RtP�ҋ�%���   �M�R`QP�҃�]� ���������������U�졀%�P���   ]��������������U�졀%�P�E���   P�҅�u]� ��%���   P�B�Ѓ�]� ��������U��E�M�UP��P�EjP�b����]��������������̸   �����������U��V�u��t���u8�EjP�b������u3�^]Ë��c����t���t��U3�;P����#�^]�����U��E��u�E�M��%��%�   ]� �����������U��E�����V��   �$�l� �   ^]á�%������%uT�EP�sW����=�.  }�����^]Ëu��t�h|�jmh�%j�G�������t ����t������%tV����x���   ^]���%    �   ^]ËM�UQR�AM������������^]�^]�K���-�%u.��L���������%��t���Fu��V� �������%    �   ^]Ã��^]Ð�� � &� z� e� � ������������U�졀%���   �BXQ�Ѓ���u]� ��%�Q|�M�RQ�MQP�҃�]� ���U�졀%���   �BXQ�Ѓ���u]� ��%�Q|�M�R8Q�MQP�҃�]� ���U��EV��j ���%�Qj j P�B�ЉF����^]� ��̡�%Vj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� ��%�Q�MP�EP�Q�JP�у��F�   ^]� ���̡�%�H���   ��U�졀%�H���   V�u�R�Ѓ��    ^]����������̡�%�P���   Q�Ѓ�������������U�졀%�P�EPQ���   �у�]� ̡�%�H�������U�졀%�H�AV�u�R�Ѓ��    ^]��������������U�졀%�H�AV�u�R�Ѓ��    ^]��������������U�졀%�P��Vh�  Q���   �E�P�ы�%���   �Q8P�ҋ�%���   ��U�R�Ѓ���^��]��������������̡�%�P�BQ�Ѓ����������������U�졀%�P�EPQ�J\�у�]� ����U�졀%�P�EP�EP�EP�EP�EPQ���   �у�]� �U�졀%�P�EP�EP�EP�EPQ�JX�у�]� �������̡�%�P�B Q��Y�U�졀%�P�EP�EP�EP�EPQ���   �у�]� �����U�졀%�P�EP�EP�EPQ�J�у�]� ������������U�졀%�H��   ]��������������U�졀%�P�R$]�����������������U�졀%�P��x  ]��������������U�졀%�P�EP�EP�EP�EPQ�J(�у�]� ��������U�졀%�P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U�졀%�P�EP�EP�EP�EPQ�J,�у�]� ��������U�졀%V��H�QWV�ҋ���%�H�QV�ҋ�%�Q�M�R4Q�MQ�MQ���W���Pj j V�҃�(_^]� �����������U�졀%�P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U�졀%�P�EP�EPQ�J@�у�]� U�졀%�P�EPQ�JD�у�]� ���̡�%�P�BLQ�Ѓ���������������̡�%�P�BLQ�Ѓ���������������̡�%�P�BPQ�Ѓ����������������U�졀%�P�EPQ�JT�у�]� ����U�졀%�P�EPQ�JT�у�]� ����U�졀%�P�EP�EPQ���   �у�]� �������������U�졀%�P�E���   ��VP�EPQ�M�Q�ҋu�    �F    ��%���   j P�BV�Ћ�%���   �
�E�P�у� ��^��]� ������̡�%�P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡�%�H�������U�졀%�H�AV�u�R�Ѓ��    ^]��������������U�졀%�P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U�졀%�P�EPQ�J�у�]� ���̡�%�P�BQ��Y�U�졀%�P�EP�EPQ�J�у�]� U��VW�������M�U�x@�EPQR���Ξ���H ���_^]� �U��VW��贞���M�U�xD�EPQR��螞���H ���_^]� �V��舞���xH u3�^�W���v����΍xH�l����H �_^�����U��V���U����xL u3�^]� W���@����M�U�xL�EPQR���*����H ���_^]� �������������U��V�������xP u���^]� W�������M�U�xP�EP�EQRP���՝���H ���_^]� ��������U��V��赝���xT u���^]� W��蟝���M�xT�EPQ��荝���H ���_^]� U���S�]��VW��t.�M��v������_����xL�E�P���Q����H ��ҍM������}��tZ��%�H�A�U�R�Ћ�%�Q�J�E�WP�ы�%�B�P�M�Q�҃���������@@��t��%�QWP�B�Ѓ�_^[��]� ������U��V���Ŝ���x` u
� }  ^]� W��譜���x`�EP��蟜���H ���_^]� ��U��VW��脜���xH�EP���v����H ���_^]� ���������U��SVW���S����x` u� }  �#���?����x`�E���P���,����H ��ҋ���%�H�]�QS�҃�;�A��%�H�QS�҃�;�,�������M�U�xD�EPQSR���؛���H ���_^[]� _^�����[]� ��������������U��V��襛���xP u
�����^]� W��荛���M�U�xP�EP�EQ�MR�UPQR���k����H ���_^]� ��������������U��V���E����xT u
�����^]� W���-����M�xT�EPQ�������H ���_^]� ��������������U��V��������xX tW�������xX�EP���ٚ���H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u��8g������t.�E�;�t'��%�J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡�%�H��   ��U�졀%�H��$  V�u�R�Ѓ��    ^]�����������U�졀%�UV��H��(  VR�Ѓ���^]� �����������U�졀%�P�EQ��,  P�у�]� �U�졀%�P�EQ��,  P�у������]� ���������̡�%�H��0  �⡀%�H��4  �⡀%�H��p  �⡀%�H��t  ��U��E��t�@�3���%�RP��8  Q�Ѓ�]� �����U�졀%�P�EPQ��<  �у�]� �U�졀%�P�EP�EP�EPQ��@  �у�]� ���������U�졀%�P�EP�EPQ��D  �у�]� �������������U�졀%�P�EPQ��H  �у�]� �U�졀%�P�E��L  ��VWPQ�M�Q�ҋu����%�H�QV�ҡ�%�H�QVW�ҡ�%�H�A�U�R�Ѓ�_��^��]� ��������������̡�%�P��T  Q�Ѓ�������������U�졀%�P�EPQ��l  �у�]� ̡�%�P��P  Q�Ѓ�������������U�졀%�P�EPQ��X  �у�]� ̡�%�H��\  ��U�졀%�H��`  V�u�R�Ѓ��    ^]�����������U�졀%�P�EP�EP�EP�EP�EPQ��d  �у�]� �U�졀%�P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���w���d����3��F�F �F$�F(�F,�F0�F4�F8�F<�F@�FD�FH�FL�FP�FT�FX�_p��G`�Gd�Gh�Gx�����G|   ��_^��������������V��W�>��t7���o����xP t$S���a���j j �XPj�FP���M����H ���[�    �~` t��%�H�V`�AR�Ѓ��F`    _^������������U��SV��Fx��%�Q��   WV�^dSP�EP�~`W�у����F|��   �> ��   �; ��   �U�~pW�^hSR��N������u#���h����%�H��0  h�   �҃��E�~P����f���j j jW�^������F|t��������F|_^[]� �F|_�Fx����^[]� �F|�����    ��%�Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��V��~d �F`tLW�};~xtBWPj�NQ��������F|u�E���~xt�    �F`_^]� �M���Fx����t�3�_^]� U��QVW�}����>+  ��%�H�QhV�҃�����%u"�H��0  h��h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���t�3�9u�~!�E���<� t��Q���)  �E��;u�|�UR�{�����_�   ^��]� �����������U��QVW�}����~*  ��%�H�QhV�҃�����%u"�H��0  h��h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���tЋE��t�3�9u�~:��E�<� t'����%�QP�Bh�Ѓ���t�M��R���,(  ��;u�|ȍEP蛘����_�   ^��]� �����������h��h�   h�%h�   �g�������t�������3��������V���(����N^�`�����������������U��VW�}�7��t��������N�`��V�M������    _^]�U��M�EV�u������t#W���    �Pf�y������f�8f�u�_^]� �U��� �E���M��"  �ȉES���V�u��W�}�ǃ��Q���ƃ��։E��B��E���؉M�E��U���M��~�U�U���)}�M��>���E��}�t�u+���I �\�P���m���u�E�����E��   )}��u��	;]��u��s���u;]�]�}�M��>P�E�V�Ѕ�}	�u���]�M��E��VP�҅��V������F��}�t!�M�+ȃ����\�P���m���u�]��;]~�����_^[��]� ���U���(W�}�����E�E���M��  �MS�؉E������ǃ��S�����E�ы���V�]�U��E܉U���]��~�E�E��)}��]��)�M�U��E�Q�M�RP������E�����E��   )}��u�;E��؉u�s���u;]�]�}�M���>P�E؋V�Ѕ�}	�u؃��]��M���E�VP�҅��i����}���F�t&�M�+ȃ���I �Pf�\����f�f�u�]��}�;E�w����%���^[_��]� ��������U���(W�}�����E�E���M��)  �ЉE������ǃ��J���SV�uƃ��ΉE��A��E����؉U��E܉M����I �U���~�M�M��)}��U��A�M�ɋE��M�t�M�+���I �\�p���m���4u�E�����E��   )}��u�;E��؉u�s���u;]�]�}�M��>P�E؋V�Ѕ�}	�u؃��]��M��E�VP�҅��Q����}���F�t�M�+ȃ���\�P������u�]��}�;E~�����^[_��]� ���������������U��E�Pu�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����E��SV��W�]�t8�u��t1�}��t*�} t$�VP��Ѕ���   |������E�   �}}_^3�[��]� �}�M���E�������uu��VP�҅�t#}����}����}��E9E�~�_^3�[��]� ��~3�E���]��]�E��E�M���؋ESP���҅�u�����_��^[��]� ���������������U����E��SV��W�]��  �u����   �}����   �} ��   �VP��Ѕ���   }�M_^�    3�[��]� �O�3����E�   �M} ����   �E���8_^3�[��]� ���M�U���<�M������uuVQ���҅�t}�O��M��W�U��M9M�~�뤅�~3�E���]��]�E��E�M���؋ESP���҅�u�����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� �����������U��V�u�F��F�����������������3  ����������D�Ez��^�P�P�]��������������N�X�N^�X]�������P�P��P(�P �P�P@�P8�P0�PX�PP�PH����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX��������U��M�A8��   �IXV�AP�I@���I�AP�I(�AX�I ���I0���A@�I �A8�I(���IH����������Dz�u�؋��5�����^��]���W���A�IX�AP�I�A8�I�A�I@�AP�I@�U��A8�IX�]������IH�����I0�����e��	����ݝx����A�I(�U��A�I �U��AX�I �]��AP�I(�����IH�E����	���������I�������]��A8�I(�A@�I �����	�������I���E��e��I0�������]��E��e����]����e��ˋE��x������]������]��AH�I@�A0�IX�����]��AX�I�AH�I(�����]��A0�I(�A@�I�����]��AP�I0�AH�I8�����]��AH�I �AP�I�����]��A8�I�A0�I �   �����]��_^��]�������U��y0 ts��U�����Au���A�Z����Au�B�Y�A�Z����Au�B�Y�A�����z��Y�A �Z����z�B�Y �A(�Z����zZ�B�Y(]� �E��Q�P�Q�P�Q �P�Q$�P�Q(�@�A,�Q�A��Q �A�A$�Q�Q(�A�A,�Q�A�A0   ]� U��y0 tL��E�A�A �A�A(�A�������������X�X�A� �A �`�A(�`�E����X�X]� ��E����������P���P�E����X�X]� ��̋�3ɉ�H�H�H�V��V�W����FP�N���3����F�F^��3���A�A�A����A�`�
�@�b�	���B�a�������U����   ��UV���q�U�W3��<��M��}���  ��S�]�k  ��؋�U��M�U��U�@�����@�U��@�B�@�������@���@�G�>��w����U���  �w������݃��B��   �U������ɋP��R�э����]��B���B�P���R���U����E������]��E��M��E������������]��E����E����E��E��]����E��]����E��]��]����U��E��U�����B���B���U������������]��E����E����������E������E��E��]����E��]����E��]����U��E��]���R�э�������B���B�P���R���U����E��������]��E����E����������E������E��E��]��E��]����E��]��U��E��]�����B���B���U����E��������]��E����E����������E������E��E��]��E��]����E��]��E��U��`�����E�U���������;���   �ލ�+���͋�@����������]��@���]��@���U������M������]��E��E����E��������]��E������������E��E��]��E��E��]����E��]��E��U�u�������������������������������M���Q�ʍU��R���[�[������E�KH��P�E��SL��H�щKP�P�ST�H�KX�P�������S\z^�E�����������zP���CP�����CX���CH���CX�������cH���[�[ �[(�C(�KP�C �KX���C�KX�C(�KH���CH�K �\���E���������za�CX�����CP�����cH�CH���CP�������[���[ �[(�CP�K(�C �KX���C�KX�CH�K(���C �KH�C�KP�����[0�[8�[@�[�CP�����CX�����KH�CX�����cP���[0�[8�[@�C8�KX�C@�KP���C@�KH�CX�K0���CP�K0�C8�KH�����[�[ �[(��$���SP������E��U�   �����}��M�����م�~�A8����u��1���U�@���K�I��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�@�K@���CX�H�D��@�����U���]��C���@�K0���CH�H���C ��C�@�K8���@�KP���C(��C�C@�H���CX�H3������U��x  �A������܃��E����E   �E�
���������ɋE������׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H�E������������������������������E����]��E��]����]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H�E��������]������M������������������������]��E��]��E��]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H���]������M������������������������]��E�Eȃ��]���E����]ȃE׃m����@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H���]������M������������������������U��E��]��E��U�������E������������;���   �P�U��+ЉU�
���������ʋE���׋��U�@���K��@�K0���CH�H���]�� �K �C�@�K8���@�KP���]�� �K(�C�C@�H���CX�H�   E)E���]����E��������������������M����������]��E��E��U�����[������_��^��]� ��[��_��^���؋�]� �����������h�%Ph_� ��������������������h�%jh_� ���������uË@����U��V�u�> t/h�%jh_� ��������t��U�M�@R�Ѓ��    ^]���U��Vh�%jh_� ���i�������t�@��t�MQ����^]� 3�^]� �������U��Vh�%jh_� ���)�������t�@��t�MQ����^]� 3�^]� �������U��Vh�%jh_� �����������t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�%jh_� ����������t�@��t�MQ����^]� 3�^]� �������U��Vh�%j h_� ���Y�������t�@ ��t�MQ����^]� 3�^]� �������U��Vh�%j$h_� ����������t�@$��t�MQ����^]� 2�^]� �������Vh�%j(h_� �����������t�@(��t��^��3�^������Vh�%j,h_� ����������t�@,��t��^��3�^������U��Vh�%j0h_� ���y�������t�@0��t�MQ����^]� 3�^]� �������U��Vh�%j4h_� ���9�������t�@4��t�M�UQR����^]� ���^]� ��Vh�%j8h_� �����������t�@8��t��^��3�^������U��Vh�%j<h_� �����������t�@<��t�MQ����^]� ��������������U��Vh�%j@h_� ����������t�@@��t�MQ����^]� ��������������U��Vh�%jDh_� ���I�������t�@D��t�MQ����^]� 3�^]� �������U��Vh�%jHh_� ���	�������t�@H��t�MQ����^]� ��������������Vh�%jLh_� �����������t�@L��t��^��3�^������Vh�%jPh_� ����������t�@P��t��^��3�^������Vh�%jTh_� ���l�������t�@T��t��^��^��������Vh�%jXh_� ���<�������t�@X��t��^��^��������Vh�%j\h_� ����������t�@\��t��^��^��������U��Vh�%j`h_� �����������t�@`��t�M�UQR����^]� 3�^]� ���U��Vh�%jdh_� ����������t�@d��t�M�UQR����^]� 3�^]� ���U��Vh�%jhh_� ���Y�������t�@h��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh�%jlh_� ���	�������t�@l��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�%jph_� ����������t�@p��t�M�UQR����^]� 3�^]� ���U��Vh�%jth_� ���y�������t�@t��t�M�UQR����^]� 3�^]� ���U��Vh�%jxh_� ���9�������t�@x��t�M�UQR����^]� 3�^]� ���U��Vh�%j|h_� �����������t�@|��t�MQ����^]� 3�^]� �������U��Vh�%h�   h_� ����������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh�%h�   h_� ���f�������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh�%h�   h_� ����������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh�%h�   h_� ����������t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U���|��A�����U����U����U��  S�V�E��EW�����������   ���������U�r�z�
�R;��4v���4��I�$ȍ��F�R�a���F�a�uB�!�]��B�a�U��B�a�U������������]��E����E����������E��������E��G��$ȍ��]��B�a�U��B�a�U������������]��E����E����������E��������E��������m�������_�U�^��[�U����U���������������������  ����������D�Ez���P�P���]� �������E�����E����X�M��X��]� �������U���@����A�������E�    ���]����]��]�����������]����]��]���   �	S�]VW�M��E����������t[��%�����E�M�����@��P������F�@��R�M������~���Q�M������v;�t�v��P�M������M����m��M�u�_^[�M�UQR�M��A�����]� ����������̋Q3���|�	��t��~�    t������u��3�������U��QV�u;��}�	���    u����;�|���^]� +ƃ�^]� �������U��VW�}��|-�1��t'�Q3���~�΍I �1�������;�t����;�|���_^]� �������������̋Q3���~%V�1�d$ ���   @u�����t������u�^�̋QV3���~�	�d$ ����Шt������u��^�������U��Q3�9A~��I ��$��������;A|�Q��~[SVW�   3ۋ���x5��%���;��E���}$��������%���;E�u�
   ���;q|݋Q���G���;�|�_^[��]�������U��	����%�����E��   @t����������wg�$�8� �E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� �� �� �� � %� ����U����S��V������   @Wt���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V��V�'v���FP�v��3����F�F^��U��SV��WV�v���^S��u���E3���;ǉ~�~t_��%�Q���   h����jIP�у�;ǉt9�}��t;��%�B���   h����    jNQ�҃����uV�u����_^3�[]� �E�~_�F^�   []� ����������U��SV��WV�Ru���^S�Iu���}3Ƀ�;��N�N��   9��   �G;���   ��%�Q���  h����jlP�у����t=� t@�G��t9��%�Jh����    ���  jqR�Ѓ����u���]���_^3�[]� �O�N�G�Q��    R�F�QP�  �����t�N�WP��QPR�h  ��_^�   []� ���������U��SV��WV�Rt���~W�It��3Ƀ�9M�N�N��   �E;���   ��    ��%�H���  h��h�   S�҃����t=�} tH�E��tA��%�Q���  h����h�   P�у����u���b���_^3�[]� �U�V�,�F   ��%�H���  h��h�   j�҃����t��E�M�F�PSPQ�a  �E����t!�V�?�W�RWP�E  ��_^�   []� ��M�_^�   []� ���U��Q2���~CS�]V�1W������������;�u��   @u�����u3���   ��
���u�_^[��]� �����������U��S�]V��3�W�~���F�F�C;CV��   �r��W�r��3��F�F��%�Q���   h��jIj�Ѓ������   ��%�Q���   h��jNj�Ѓ����uV�Fr����_��^[]� ��F   �F   ����K�H�C��B�_��^�   []� � r��W��q��3��F�F��%�B���   h��jIj�у����t[��%�B���   h��jNj�у�����\�����F   �F   ����S�Q��K�H��C�B��   _��^[]� �����������U��3�V���F�F�F�EP�������^]� �������������U��EVP���������^]� ����������U��U��t�M��t�E��tPRQ�   ��]������������V��F��Wu�~��N�ɍ<u�< ��u_3�^á�%�H�F��  h<�j8��    RP�у���tщ~�F_�   ^���U��V��F;Fu������u^]� �N�V�E���   F^]� �����������U��V��FW�};�~ ��|�F�M��_�   ^]� _3�^]� })�V;Vu��������t�F�N��    �F9~|׋V;Vu���������t��F�N�U���F_�   ^]� ������U��V��FW�};�~����}3�;Fu������u_^]� �F;�~�N�T������;ǉ�F�M���F_�   ^]� �U��E��|4�Q;�}-���;Q}V�d$ �Q�t������2;A|�^�   ]� 3�]� ������������U��Q3���V~�I�u91t����;�|���^]� �������V��W�~W��n��3����_�F�F^�����A    ��������̋Q�B���|;�}�QV�4���tP�1�����^�3�����������̍Q3��Q�Q�A�Q�A������������W���O�G;�t#��tV�q��t�~ u3���j�҅���u�^�G�G�G�G    �G�G    _�����U��A��3�;�Vt!��t�M���;�t�@��t
�x t��u�3�^]� ��������U��Q�E�P�Q�P�Q�B�A]� �U��E�Q�P�Q�P�Q�B�A]� ̋Q��3�;�t�ʅ�t�I����t
�y t��u�����������U��E�P�Q�H�A�@�H]� ����U��E�P�Q�H�A�A�H]� ���̋Q��t!�A��t�B�A�Q�P�A    �A    ��������V��W�~W�|���l��3����_�F�F^��������������U���SV�uW���^S�}��l��3���F�F�O�N�W���V9G�E~��I �O���F9F�U�uL��u�~��~��t���< ��t\��%�H���  h<�j8��    RP�у���t3�~�}���V��M����E�F��;G�E|�_^�   [��]� _^3�[��]� �������������U��V�u��|'�A;�} �U��|;�};�t�A��W�<��<���_^]� ���������U��EV�u;�}����|,�Q;�}%��|!;�};�t�QW�<�P������tVW����_^]� ����������U��V�q3���W~�Q�}9:t����;�|���P�����_^]� ���������������U����E�Qj�E��ARP�M��E����������]� �����U����Q�Ej�E��A�MRPQ�M��E���������]� ̋A��;�t?W3�;�t7V�H;�t	9yt���3��P;�t;�t�J�H�P�Q�x�x;���u�^_������̋Q���8�t!�A��t�B�A�Q�P�A    �A    �̋�� ���@8��HV3��q�q�P�r�r�8��p�p�p�P�H^������V����������F3�;��F8�t�N;�t�H�F�N�H�V�V�F;��F8�t�N;�t�H�F�N�H�V�V^�U��E�UP�AR�Ѓ�]� ���������U��V��N3�;��8�t�F;�t�A�F�N�H�V�V�Et	V�fl������^]� ������������U��V��W�~W�|���h��3����E��F�Ft	V�!l����_��^]� ������U��V��������Et	V��k������^]� ��������������̋T$�L$��ti3��D$��u��   r�=�A t�  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$øS!����O����A�������� �����7���������  �|$ ��%t�.  ���Q����  Y�V��������D$tV��j��Y��^� U��Q�E��SVW�  ����   Wj ��P������u3��  V�>����Vj u��P���ދF�~�E�F�E�F�E����  ��P���E��t�� �  �M���%�E�����j��%��%��%�=�%�z)  ��Y�s����q  ��u
�)  �`����(  ����A�q'  ��%�!  ��}�&  ���&  ��| �"$  ��|j �  ��Yu��%�   �#  ��3�;�u59=�%�������%9=(&u��  9}u{�#  ��  �%)  �j��uY�}  h  j�|   ��;�YY�����V�5�58&��  Y�Ѕ�tWV�  YY� ��N���V�  Y�m�����uW��  Y3�@_^[�� jh��*  ����]3�@�E��u9�%��   �e� ;�t��u.�����tWVS�ЉE�}� ��   WVS������E����   WVS�Y����E��u$��u WPS�E���Wj S���������tWj S�Ѕ�t��u&WVS�~�����u!E�}� t�����tWVS�ЉE��E������E���E��	PQ�)  YYËe��E�����3���)  Ã|$u�+  �t$�L$�T$�����Y� ;�u����,  QSUVW�5�A�f  �5�A���t$�U  ��;�YY��   ��+ލk��rxV�-  ��;�YsJ�   ;�s���;�rP�t$��  ��YYu�F;�rCP�t$��  ��YYt3��P�<��u  Y��A�t$�f  ���W�[  Y��A�D$Y�3�_^][Y�Vjj �5  ��V�4  ������A��AujX^Ã& 3�^�jh��(  ��  �e� �u�����Y�E��E������	   �E��(  ���  ��t$���������YH�jh �5(  �e� �u;5�@w"j�.  Y�e� V��6  Y�E��E������	   �E��A(  �j�-  Y�U�l$�����   S��VW3�95T'��u�;  j�n9  h�   �#  YY��@��u;�t���3�@P���uU�S���;�Yu;�u3�G�����WV�5T'�Ӌ���u&9�.j_tU�n;  ��Yu���;  �8�;  �8_��^[]�U�L;  Y��:  �    3�]�jh �#'  �u��tu�=�@uCj�-  Y�e� V��-  Y�E��t	VP�.  YY�E������   �}� u7�u�
j�u,  Y�Vj �5T'����u�w:  ����P�.:  �Y��&  ���������̃=�A t-U�������$�,$�Ã=�A t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$�������U��WV�u�M�}�����;�v;���  ��   r�=�A tWV����;�^_u^_]�T;  ��   u������r*��$����Ǻ   ��r����$���$����$�(���#ъ��F�G�F���G������r���$���I #ъ��F���G������r���$���#ъ���������r���$���I �xph`XPH�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$���������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�0�����$���I �Ǻ   ��r��+��$�4�$�0�Dh��F#шG��������r�����$�0�I �F#шG�F���G������r�����$�0��F#шG�F�G�F���G�������V�������$�0�I ����'�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�0��@HXl�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̃��$�;  �   ��ÍT$�h;  R��<$�D$tQf�<$t� ;  �   �u���=�% ��;  �   ���;  �  �u,��� u%�|$ u����:  �"��� u�|$ u�%   �t����-@�   �=�% �6;  �   ���?:  Z�U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]Ã%�A �p;  ��A3�ËD$��V���F uc��  �F�Hl��Hh�N�;xt���Hpu�E  ��F;�t�F���Hpu�=  �F�F�@pu�Hp�F�
���@�F��^� U���V�u�M��l����u�P��G  ��e�F�P�F  ��Yu��P��G  ��xYuFF�M����   �	��	�F�����F��u�8M�^t�E��`p���U���V�u�M�������E��ɋu�t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B�Ɉu��}� ^t�E��`p�����D$�����Az3�@�3��U��QQ�} �u�ut�E�P�	G  �M��E��M��H��EP�G  �E�M�����j �t$�t$�t$������Å�V��tV�K  @PV�V�H  ��^�j �t$�z���YY�j �t$�����YY�U���SVW�u�M��������3�;�u+�I2  j_VVVVV�8�D  ���}� t�E��`p����!  9uv�9u~�E�3���	9Ew	�2  j"뺀} t�U3�9u��3Ƀ:-����ˋ��:����}�?-��u�-�s�} ~�F�����E����   � � �3�8E��E��}�u����+�]h��SV��J  ��3ۅ�tSSSSS��B  ��9]�Nt�E�GF�80t.�GHy���-F��d|
�jd_�� ��F��
|
�j
_�� �� F�D/t�90uj�APQ�F  ���}� t�E��`p�3�_^[��U���,��3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�L  3ۃ�;�u��0  SSSSS�0�C  �����o�E;�v����uu����3Ƀ}�-��+�3�;���+��M�Q�NQP3��}�-��3�;�����Q�;J  ��;�t���u�E�SP�u��V�u��������M�_^3�[�������U��j �u�u�u�u�u������]�U���$VW�u�M��E��  3��E�0   �k���9}}�}�u;�u+��/  j^WWWWW�0�B  ���}� t�E�`p����  9}vЋE��9E� w	�/  j"���}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW� �������t�}� � ��  �M�ap��  �;-u�-F�0F�} je����$�x�FV�c6  ��YY�L  �} ���ɀ����p��@ �2  %   �3��t�-F�]�0F������$�x��OF��ۃ����  �3���'3��u!�0�O����� F�u�U���E��  ��1F��F9U�Eu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~M�W#U���M�#E���� ��J  f0 ��f=9 vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �J  f= v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V�/�����u�E�8 u���} �4����$�p���WF�#J  3�%�  #�+E�SY�x;�r�+F�
�-F�����;Ӌ��0|$��  ;�rSQRP��H  0�F;��U�����u��|��drj jdRP��H  0��U�F����;�u��|��
rj j
RP�H  0��U�F���]�0��F �}� t�E�`p�3�[_^��U���SVW�u�؋s���M�N������u-�{,  j^�03�PPPPP�>  ���}� t�E��`p����   �} v̀} t;uu3��;-����� 0�@ �;-��u�-�w�C3�G�����n����0F���} ~D���Y����E����   � � ��[F��}&�ۀ} u9]|�]�}���(���Wj0V�k������}� t�E��`p�3�_^[��U���,��3ŉE��ESVW�}j^V�M�Q�M�Q�p�0��F  3ۃ�;�u�n+  SSSSS�0�=  �����Z�E;�v���u��3Ƀ}�-��+��u�M�Q�M��QP3��}�-���P��D  ��;�t���u�E�SV�u���d������M�_^3�[������U���0��3ŉE��ESV�uWj_W�M�Q�M�Q�p�0�F  3ۃ�;�u�*  SSSSS�8��<  �����   �M;�vދE�H�E�3��}�-������<0u��+ȍE�P�uQW�ED  ��;�t��X�E�H9E������|-;E}(:�t
�G��u��_��u�E�j�u���u��������u�E�jP�u���u�u�������M�_^3�[������U��E��et_��EtZ��fu�u �u�u�u�u�&�����]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u������u �u�u�u�u�u�|�����]�U��j �u�u�u�u�u�u�^�����]�VW3�����6�  ����(Y�r�_^�Vh   h   3�V�F  ����tVVVVV�c:  ��^�U�������]�����]��E��u��M��m��]����]�����z3�@��3���h��� ���th��P����tj �������jh@��  j�O  Y�e� �u�N��t/��%��%�E��t9u,�H�JP�u���Y�v�l���Y�f �E������
   ��  Ë���j�  Y���������������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t�����&'  �t$�}%  �5��  h�   �Ѓ��h��� ���th��P����t�t$����t$�����Y�t$�$��j��  Y�j�  Y�V������t�Ѓ�;t$r�^�V�t$3����u���t�у�;t$r�^ËL$V3�;�u��&  VVVVV�    �%9  ��jX^á�%;�tډ3�^ËD$V3�;�u�&  VVVVV�    ��8  ��jX^�95�%tۋ�%�3�^Ã=�� th���YD  ��Yt�t$���Y����hD�h,��6�����YYuTVWhA4�(���� ��ƿ(�;�Ys���t�Ѓ�;�r�=�A _^th�A��C  ��Ytj jj ��A3��jh`�&  j�  Y3��}�3�C9,&t~�(&�E�$&9}u[�5�A��  �E��5�A��  YY���u�9}�t&���u�;u�r�> t��>�  ;�t�W�  Y����hT��H��2���Yh\��X��"���Y�E������   �} u(�,&j�  Y�u�����3�C�} tj��  Y��  �j j�t$�������jj j �������V�   ��V�%%  V��E  V�6  V�2&  V��E  V�C  V�  V�C  h�%�v   ��$�^�U��QQSV3��E�F3�P�u��]�������}�Y~���BWS� ��p<�f9^�F�|0v#Wh��0�����YYt�FC��(;�r���e� �E�_^[��V�5�5(��օ�t!����tP�5���Ѕ�t���  �&h�� �����t#�J�����th�V����t
�t$�ЉD$�D$^�j ����Y�V�5�5(��օ�t!����tP�5���Ѕ�t���  �&h�� �����t#�������th,�V����t
�t$�ЉD$�D$^��,�� V�5�(�����u�54&�k���Y��V�5�0���^á���tP�5<&�A���Y�Ѓ�����tP�4����i  jh��  h�� ��E�u�F\h3�G�~��t/������t&h��u���Ӊ��  h,��u��Ӊ��  �~pƆ�   CƆK  C�p�FhP�8�j�  Y�e� �E�Fl��u�x�Fl�vl�1  Y�E������   �  �j�  Y�VW���5�������Ћ���uNh  j�  ����YYt:V�5�58&����Y�Ѕ�tj V�����YY� ��N���	V�����Y3�W�<�_��^�V��������uj�����Y��^�jh���  �u����   �F$��tP�z���Y�F,��tP�l���Y�F4��tP�^���Y�F<��tP�P���Y�FD��tP�B���Y�FH��tP�4���Y�F\=htP�#���Yj��  Y�e� �~h��tW�@���u��ptW�����Y�E������W   j�  Y�E�   �~l��t#W��0  Y;=xt���t�? uW��.  Y�E������   V����Y�  � �uj�]  YËuj�Q  YÃ=�tLW�|$��u&V�5�5(��օ�t�5�5���Ћ�^j �5�58&�`���Y��W����_����t	j P�0��Wh�� �����u	�����3�_�V�5�h\�W��hP�W�0&��hD�W�4&��h<�W�8&�փ=0& �50��<&t�=4& t�=8& t��u$�(��4&�4��0&u'�58&�<&�,�������   �54&P�օ���   �J����50&������54&�0&������58&�4&������5<&�8&��������<&�7  ��teh;)�50&����Y�Ѓ���tHh  j�   ����YYt4V�5�58&�����Y�Ѕ�tj V�����YY� ��N��3�@��l���3�^_�VW3��t$���������Yu'9@&vV�D����  ;@&v��������uɋ�_^�VW3�j �t$�t$�@  ������u'9@&vV�D����  ;@&v��������u���_^�VW3��t$�t$��@  ����YYu-9D$t'9@&vV�D����  ;@&v��������u���_^�jTh���	  3��}��E�P�T��E�����j@j ^V�@���YY;��  ��@�5�@��   �0�@ ���@
�x�@$ �@%
�@&
�x8�@4 ��@��@��   ;�r�f9}��
  �E�;���   �8�X�;�E�   ;�|���E�   �[j@j ����YY��tV�M����@���@ ��   �*�@ ���@
�` �`$��@%
�@&
�`8 �@4 ��@��;�r��E�9=�@|���=�@�e� ��~m�E����tV���tQ��tK�uQ�P���t<�u���������4��@�E� ���Fh�  �FP�O=  YY����   �F�E�C�E�9}�|�3ۋ���5�@����t���t�N��r�F���uj�X�
��H������P�L������tC��t?W�P���t4�>%�   ��u�N@�	��u�Nh�  �FP�<  YY��t7�F�
�N@�����C���g����5�@�H�3��3�@Ëe��E����������  �VW��@�>��t1��   �� t
�GP�X����@   ;�r��6�/����& Y�����A|�_^�S3�9�AVWu�)  �5�%3�;�u����   <=tGV��3  Y�t�:�u�jGW������;�YY�=&tˋ5�%U�@V�3  ��E�>=Yt/jU�Z���;�YY�tJVUP��3  ����tSSSSS��+  �����8u��5�%�r�����%���A   3�Y]_^[��5&�M����&�����U��Q�MS3�9EV���U�   t	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�C?  ��Yt��} t
�M��E�F�ۋU�Mt2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=����Pt#�^>  ��Yt��M�E�F��M��E���;>  ��YtF���UF�V�����t� B�U��M�����E��^[t�  ���U���S3�9�AVWu�&  h  �H&VS�L'�\���A;É5&t8�E�u�u��U��E�PSS�}������E���=���?sJ�M���sB�����;�r6P������;�Yt)�U��E�P�WV�}�������E���H� &�5&3�����_^[��QQ�P'SUVW�=p�3�3�;�j]u-�׋�;�t�P'   �"����xu	�ţP'��P'����   ;�u�׋�;�u3���   f9��t�f9u��f9u�=l�SSS+�S��@PVSS�D$4�׋�;�t2U�����;�Y�D$t#SSUP�t$$VSS�ׅ�u�t$�/���Y�\$�\$V�h����X;�t;�u��d���;��p���8t
@8u�@8u�+�@��U�Z�����;�YuV�`��D���UVW������V�`���_^][YY�VW����;ǋ�s���t�Ѓ�;�r�_^�VW����;ǋ�s���t�Ѓ�;�r�_^�U��QQV�E�3�P�u��u��U�����YtVVVVV�'  ���E�P�q�����YtVVVVV�t'  ���}�^u�}�r3�@��jX��3�9D$j ��h   P�x����T'u3���}�������@u$h�  �  ��Yu�5T'�t��%T' ��3�@�U3�=�@uTS��W3�9-�@~1V�5�@��h �  U�v��|��6U�5T'�Ӄ�G;=�@|�^�5�@U�5T'��_[�5T'�t��-T']��U��QQV���������F  �V\��W�}��S99t��k����;�r�k��;�s99u���3���t
�X�ۉ]�u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   ���=����;�}$k��~\�d9 �=���B߃�;�|�]�� =�  ��~du	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�øcsm�9D$u�t$P����YY�3��hp7d�5    �D$�l$�l$+�SVW��1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q���������������̃�S�\$ UV�s35�W�����D$ �D$   �{t�N�38������N�F�38������D$(�@f�  �k����L$0�T$�D$�L$ �S�t^�Dm �L��ɍ\���D$t���<9  ���D$|DL�D$�����ù|$ t$����t�N�38�S����N�F�38�C����D$_^][����D$    �ƋL$(�9csm�u*�=�@ t!h�@�<0  ����t�T$(jR��@���L$,��8  �D$,9hth�W�Ջ���8  �D$,�L$�H����t�N�38�����N�V�3:�����K���l8  �{��P���h�W�˺�����8  ����U������e� �e� SW�N�@�;ǻ  ��t��t	�У��`V�E�P����u�3u����3�� �3����3��E�P����E�3E�3�;�u�O�@����u������5��։5�^_[��U��� S3�9]u �  SSSSS�    �Y#  ������   �M;�V�ut!;�u��  SSSSS�    �*#  ������S����;ȉE�w�M�W�u�E��u�E�B   �u�u�P�u��y9  ��;��t�M�x�E����E�PS�Y7  YY��_^[���t$j �t$�t$�t$�8������U���(  �`(�\(�X(�T(�5P(�=L(f�x(f�l(f�H(f�D(f�%@(f�-<(��p(�E �d(�E�h(�E�t(��������'  �h(�d'�X'	 ��\'   ���������������������'j��A  Yj ���hh�����=�' uj��A  Yh	 ����P�����jh�����3��]3�;���;�u�<  �    WWWWW�{!  ������S�=�@u8j��  Y�}�S�?  Y�E�;�t�s���	�u���u��E������%   9}�uSW�5T'��������R����3��]�u�j�   Y�VW3���*�<��u����8h�  �0���/  ��YYtF��$|�3�@_^Ã$�� 3���S�X�V��W�>��t�~tW��W�`����& Y����|ܾ�_���t	�~uP�Ӄ���|�^[�U��E�4�����]�jh�<���3�G�}�3�9T'u�r  j��  h�   ����YY�u�4��9t���nj�<���Y��;�u�  �    3��Qj
�Y   Y�]�9u,h�  W�.  YY��uW����Y�x  �    �]���>�W�u���Y�E������	   �E�������j
�*���Y�U��EV�4���> uP�$�����Yuj����Y�6���^]�h@  j �5T'������@uËL$�%�+ �%�@ ��@3���@��@   @Ë�@��@k����T$+P��   r	��;�r�3��U����M�AV�uW��+y�������i�  ��D  �M��I���M���  S�1��U�V��U��U����]ut��J��?vj?Z�K;KuB�� �   �s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J;։M�v��;�t^�M�q;qu;�� �   �s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���� �Ls%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   ��+����   ��@�5|�h @  ��H� �  SQ�֋�@��+�   ���	P��+�@��@����    ��+�@�HC��+�H�yC u	�`���+�x�ueSj �p�֡�+�pj �5T'����@��+k���@+ȍL�Q�HQP�:  �E����@;�+v�m��@��@�E��+�=�@[_^�á�@V�5�@W3�;�u4��k�P�5�@W�5T'���;�u3��x��@�5�@��@k�5�@h�A  j�5T'��;ǉFt�jh    h   W���;ǉFu�vW�5T'��뛃N��>�~��@�F����_^�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W�����u����   �� p  ;��U�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[��U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I��?�M�vj?Y�M��_;_uC�� �   �s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O��?�L1�vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���� �Ls�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N��?�]�K�vj?^�E���   �u���N��?vj?^�O;OuB�� �   �s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���� �Ls�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[��U�����@�Mk��@������M���SI�� VW}�����M���������3���U���@����S�;#U�#��u
��;؉]r�;�u��@��S�;#U�#��u
��;ى]r�;�u[��{ u
���];�r�;�u1��@�	�{ u
��;ى]r�;�u�����؅ۉ]u3��	  S�@���Y�K��C�8�t��@�C�����U�t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��ɍy�>u;�+u�M�;�@u�%�+ �M���B_^[��QS�\$VW3�3�;�tG��r���w  Uj�:7  ��Y�1  j�)7  ��Yu�=�%�  ���   �?  h��  S��+U�  ����tVVVVV��  ��h  ��+Vj ��, �\���u&h �h�  V��  ����t3�PPPPP�  ��V�.  @��<Yv8V�!  ��;�j��.h��+�QP�5  ����t3�VVVVV�^  ���3�h��SU�&5  ����tVVVVV�:  ���4�SU�5  ����tVVVVV�  ��h  h��U�#3  ���3j��L���;�t%���t j �D$P�4��6�n  YP�6U���]_^[Y�j�5  ��Ytj�5  ��Yu�=�%uh�   �4���h�   �*���YYËD$3�;��tA��-r�H��wjXË���D���jY;��#�����������u�0Ã���������u�4Ã��V������L$Q�����Y��������0^ËD$��.��5�.�������Yt�t$�Ѕ�Yt3�@�3��U��$X�����(  ��3ŉ��  �8Vtj
�P���Y�  ��tj�  Y�8��   ���   ���   ���   �]|�ux�}tf���   f���   f�]pf�Elf�ehf�md����   ���  ���  ���   �E�  ���   �@�jP���   �E�j P�y����E����EЍE�j �E�  @�u��E�����E�P���j����̋D$��.�U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]��̀zuf��\���������?�f�?f��^���٭^����\�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^����\�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp����T���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-@��p��� ƅp���
��
�t���������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR��0  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   ��@��   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z��l������������\������   s��|���d������������T������   v��t��jh(�����e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E������U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�^�����t3�@�3�[��������A3���������U��W�}3�������ك��E���8t3�����_��-�  t"��t��tHt3�ø  ø  ø  ø  �SUVW�  ��U3��^WS�ܶ���~�~�~3��~����p��+Ɗ�CMu���  �   ��ANu�_^][�U��$d�����  ��3ŉ��  SW�E�P�v������   ��   3����  @;�r�E���ƅ�   t+�]����;�w+�@P���  j R�,�����C�C��u�j �v�E��vPW���  Pjj �3  3�S�v���  WPW���  PW�vS�1  ��DS�v���  WPW���  Ph   �vS�g1  ��$3��LE���t�L���  ���t�L ���  ��  �Ƅ   @;�r��M��  �E�����3�)E��U���  ЍZ ��w�L�р� ���w�L �р� ���  A;�rŋ��  _3�[�/����Ŝ  ��jhH�������������Gpt�l t�wh��uj ����Y�������j�����Y�e� �wh�u�;5�t6��tV�@���u��ptV����Y���Gh�5��u�V�8��E������   뎋u�j����Y�U���S3�S�M��3������� /u� /   ���8]�tE�M��ap��<���u� /   ����ۃ��u�E��@� /   ��8]�t�E��`p���[��U��� ��3ŉE�S�]V�uW�h�����3�;��}u�������3��  �u�3�9����   �E��0=�   r����  �f  ����  �Z  ��P������H  �E�PW������)  h  �CVP�V���3�B��9U�{�s��   �}� ��   �u�����   �F����   h  �CVP�����M��k�0�u�����u��*�F��t(�>����E����D;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   ����j�C�C���Zf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�.����C�S��s3��{����95 /�b�������M�_^3�[�2�����jhh�����M���������}�������_h�u�����E;C�W  h   ����Y�؅��F  ��   �wh���# S�u�����YY�E�����   �u��vh�@���u�Fh=ptP�����Y�^hS�=8����Fp��   ����   j�v���Y�e� �C�/�C�/�C�/3��E��}f�LCf�E/@��3��E�=  }�L���@��3��E�=   }��  ���@���5��@���u��=ptP�>���Y��S���E������   �0j�����Y��%���u ��ptS����Y������    ��e� �E��b���Ã=�A uj��V���Y��A   3��SUV�t$���   3�;�Wto=`th���   ;�t^9(uZ���   ;�t9(uP蒶�����   ��/  YY���   ;�t9(uP�q������   �p/  YY���   �Y������   �N���YY���   ;�tD9(u@���   -�   P�-������   ��   +�P�������   +�P�������   ���������   �=�t9��   uP�[-  �7�ڵ��YYj�~P[���t�;�t9(uP蹵��Y9o�t�G;�t9(uP袵��Y��Ku�V蕵��Y_^][�SUV�t$W�=8�V�׋��   ��tP�׋��   ��tP�׋��   ��tP�׋��   ��tP��j�^P]�{��t	���tP�׃{� t
�C��tP�׃�Mu؋��   �   P��_^][�V�t$��tSUW�=@�V�׋��   ��tP�׋��   ��tP�׋��   ��tP�׋��   ��tP��j�^P]�{��t	���tP�׃{� t
�C��tP�׃�Mu؋��   �   P��_][��^Å�t7��t3V�0;�t(W�8�������YtV�R����> Yu���tV�x���Y��^�3��jh��b����x������Fpt"�~l t�a����pl��uj �X���Y���u����j����Y�e� �Fl�=x�i����E��E������   ��j����Y�u�ËD$�@/�U��$X�����(  ��3ŉ��  V���   ���   ���   �]|�ux�}tf���   f���   f�]pf�Elf�ehf�md����   ���  ���  ���   �E�  ���   �@�jP���   �E�j P�Ŭ���E��EЍE؃��E�  ��u��E����j ������E�P�����u��uj�C   Yh  ����P������  3�^�t����Ũ  ��U���5@/�������Yt]��j��  Y]�����U����u�M�������E����   ~�E�Pj�u��,  ������   �M�H���}� t�M��ap��Ã=/ u�D$�h�A���j �t$����YY�U���SV�u�M������]�   ;�sT�M胹�   ~�E�PjS�W,  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�,  ��YYt�Ej�E��]��E� Y��`���� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�&  ��$���o�����u�E���M�3��e���}� t�M��ap�^[�Ã=/ u�D$�H���w�� �j �t$�����YY�U���(��3ŉE�SV�uW�u�}�M��0����E�P3�SSSSW�E�P�E�P�6  �E�E�VP�,  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[������U���(��3ŉE�SV�uW�u�}�M�芶���E�P3�SSSSW�E�P�E�P��5  �E�E�VP�0  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�H���������U��WV�u�M�}�����;�v;���  ��   r�=�A tWV����;�^_u^_]�4�����   u������r*��$��a��Ǻ   ��r����$��`�$��a��$�Ha��`a(a#ъ��F�G�F���G������r���$��a�I #ъ��F���G������r���$��a�#ъ���������r���$��a�I �a�a�a�a�axapaha�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��a���a�a�a�a�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�Pc�����$� c�I �Ǻ   ��r��+��$�Tb�$�Pc�db�b�b�F#шG��������r�����$�Pc�I �F#шG�F���G������r�����$�Pc��F#шG�F�G�F���G�������V�������$�Pc�I cccc$c,c4cGc�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�Pc��`chcxc�c�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�ËL$S3�;�VWt�|$;�w�r���j^�0SSSSS���������1�t$;�u��ًъ�BF:�tOu�;�u��6���j"Y�����3�_^[�U��MSV�u3�;�W�yu����j^�0SSSSS�M��������   9]v݋U;ӈ~���3�@9Ew�����j"Y�����;��0�F~�:�t��G�j0Y�@J;��M;ӈ|�?5|�� 0H�89t�� �>1u�A��~W�f���@PWV�������3�_^[]�U��Q�U�BS��VW��% �  ��  #ωE�B��پ   �%�� �ۉu�t;�t�� <  �(��  �$3�;�u;�u�Ef�M�X��L��<  �]����������M��E���ΉH�u��P������Ɂ���  �։P�t�M�_^f�H[��U���0��3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���u�����f��"6  �uЉC�E։�EԉC�E�P�uV������$��t3�PPPPP�������M�_�s^��3�[�ަ��������������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j�r���Y�U��E�M%����#�������Vt1W�}3�;�tVV�>  YY������j_VVVVV�8��������_��u��P�ut	�`>  ���W>  YY3�^]��������������̋L$f�9MZt3�ËA<��8PE  u�3�f�x�����������̋D$�H<��ASV�q3҅�W�Dv�|$�H;�r	�X�;�r����(;�r�3�_^[���������������U��j�h�hp7d�    P��SVW��1E�3�P�E�d�    �e��E�    h   �<�������tU�E-   Ph   �R�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]�jh�����觿���@x��t�e� ���3�@Ëe��E��������������hki����Y��/ËD$��/��/��/��/ËD$��V9Pt��k�t$��;�r�k�L$^;�s9Pt3���5�/�����Y�j h������3��}�}؋]��Lt��jY+�t"+�t+�td+�uD�e������}؅�u����a  ��/��/�`�w\���`���������Z�Ã�t<��t+Ht�<����    3�PPPPP�y�����뮾�/��/���/��/�
��/��/�E�   P�6����E�Y3��}���   9E�uj�˺��9E�tP����Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.���M܋����9M�}�M�k��W\�D�E���螻����E������   ��u�wdS�U�Y��]�}؃}� tj ����Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3�����ËD$��/ËD$��/��t$���3�@� jh����3��}��5�/����Y��;�uS�E�P�·��Y;�tWWWWW��������}�t!hP�� �;�th(�P����;�u��kV�=���Y��/�}��u�u�։E��/�E� � �E�3�=  �����Ëe�}�  �uj�<��e� �E������E������jh(�T����M3�;�v.j�X3���;E�@u������    WWWWW�5�����3���   �M��u;�u3�F3ۉ]���wi�=�@uK������u�E;�@w7j�Z���Y�}��u����Y�E��E������_   �]�;�t�uWS������;�uaVj�5T'����;�uL9=�.t3V����Y���r����E;��P����    �E���3��uj� ���Y�;�u�E;�t�    �������jhH�6����]��u�u�5���Y��  �u��uS����Y�  �=�@��  3��}�����  j�g���Y�}�S�����Y�E�;���   ;5�@wIVSP��������t�]��5V�|���Y�E�;�t'�C�H;�r��PS�u�谢��S�����E�SP������9}�uH;�u3�F�u������uVW�5T'���E�;�t �C�H;�r��PS�u��\���S�u��Z������E������.   �}� u1��uF������uVSj �5T'�������u�]j����YË}����   9=�.t,V�����Y�����������9}�ul����P�?���Y��_����   �h���9}�th�    �q��uFVSj �5T'�������uV9�.t4V����Y��t���v�V�p���Y�����    3�������	����|�����u���������P�����Y����U����u�M��R����E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap���jj �t$j ����������SVW�T$�D$�L$URPQQh�pd�5    ��3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C��:  �   �C��:  �d�    ��_^[ËL$�A   �   t3�D$�H3�芜��U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�:  3�3�3�3�3���U��SVWj j hqQ��^  _^[]�U�l$RQ�t$������]� U��QV�uV��D  �E�F��Yu����� 	   �N ����-  �@t������ "   ��S3ۨt��^��   �N�����F�F����f��F�^�]�u,��B  �� ;�t�B  ��@;�u�u�LB  ��YuV��A  Yf�FW��   �F�>�H��N+�I;��N~WP�u��@  ���E��M�� �F����y�M���t���t������������@�� �@ tjSSQ�l9  #����t%�F�M��3�GW�EP�u�@  ���E�9}�t	�N �����E%�   _[^���A@t�y t$�Ix��������QP�z���YY���u	���U��V����M�E�M�����>�t�} �^]��G@SV����t4� u.�D$�-��L$������C�>�u�C����8*u�ϰ?�i����|$ �^[�U��$�����x  ��3ŉ��  ��   S��  V3�W��  ��  �M��EЉ}ԉu��u�u��u��uĉu��u��M���9u�u-�����VVVV�    V�������}� t�E��`p������  �E��@@��   P�@B  ���Yt6�u��2B  ���Yt(�u��$B  �u����4��@�B  ����YY3��� �@$�u����u���A  ���Yt6�u���A  ���Yt(�u���A  �u����4��@�A  ����YY3��� �@$��"���;������3Ʉ҉ủu؉u��U���  C�}� �]���  ��, <Xw����X���3��3�3����x�j��Y;��E��z  �$�}�M���u��u��u��uĉu�u��X  �� t>��t-��tHHt���9  �M��0  �M��'  �M��  �M�   �  �M��	  ��*u ���}ԋ�;��}���  �M��]���  �E�k�
�ʍDЉE���  �u���  ��*u���}ԋ�;��}���  �M���  �E�k�
�ʍDЉE��  ��ItF��ht8��lt��w�x  �M�   �l  �;luC�M�   �]��W  �M��N  �M� �E  �<6u�{4uCC�M� �  �]��(  <3u�{2uCC�e�����]��  <d�  <i��  <o��  <u��  <x��  <X��  �u��E�P��P�u��  Y���E�Yt�MЍu�������C���]���  �MЍu�������  ��d�r  ��  ��S��   tZ��AtHHt@HHtHH�N  �� �E�   �U�M�@9u��]�   �]܉E���  �E�   �	  f�E�0uu�M�   �lf�E�0u�M�   �M����u������f�E��}ԋ��}���  ;�u���E܋E��E�   �  ��X�9  HHt]+��d���HH��  ��f�E��}�t'�G�Ph   �E�P�E�P��?  ����t�E�   ��G��E��E�   �E�E��P  ���;Ɖ}�t.�H;�t'f�E� � �M�t�+����E�   �  �u��  ���E�P����Y��  ��p��  �t  ��e��  ��g�������itY��nt��o��  �E��E�   tI�M�   �@�7���}��=  ����  �E� t	f�E�f���Ẻ�E�   �  �M�@�E�
   �M�f���C  ��W���k  u��guG�E�   �>9E�~�E��}�   ~-�u���]  V�ز�����U�Y�E�t
�E܉u�����E�   3�����E��G��E��E�P�u����u��}�P�u��E�SP�5��F���Y�Ћ}����   t9u�u�E�PS�5�� ���Y��YY�}�gu;�u�E�PS�5�����Y��YY�;-u�M�   C�]�S�r����E�   �M��!��s�p���HH��������Y  �E�'   �E��E�   ������E�Q�E�0�E��E�   ����f�� ��������� t��@�}�t�G���G�����@�G�t��3҉}���@t;�|;�s�؃� �ځM�   f�E� ��ڋ�u3ۃ}� }	�E�   ��e���   9E�~�E����u!Eč��  �E��M������t$�EؙRPSW�Z.  ��0��9�]�����~M��N�̍��  +�Ff�E� �E؉u�tL��t�΀90tA�M܋M��0@�2If90t@@;�u�+E����;�u���E܋E��I�8 t@;�u�+E܉E؃}� ��   �E�@t%f� t�E�-��t�E�+��t�E� �E�   �]�+]�+]��E�u�uЍE�Sj �;������uċ}ЍE̍M��K����E�Yt�E�uWSj0�E��������}� �E�tQ��~M�u܉E���M�Pj���  P�E�FPF��;  ����u9E�t�u��E̍��  ������}� Yu���M����M�P�E������Y�}� |�E�tWSj �E��������}� t�u��&����e� Y�]�����E�t$�M��}Ԋ��)���������    3�PPPPP�$����}� t�E��`p��E̋��  _^3�[�z������  ���vEu`u�u�u�u(v w�%�@ �U��� SVW踩��3�9�/�E��]��]�]���   h8������;��y  �5�h,�W��;��c  P������$�W��/��P�����$�W��/��P�ը����/�E�P������YYtSSSSS�A������}�u,h��W��P蠨��;�Y��/th��W��P舨��Y��/��/�M�;�ty9�/tqP�ߨ���5�/���Ҩ��;�YY��tV;�tR��;�t�M�Qj�M�QjP�ׅ�t�E�u3�E�P蟥����YtSSSSS�������}�r	�M    �D�M   �;��/;E�t1P�d���;�Yt&��;ÉE�t��/;E�tP�F���;�Yt�u��ЉE��5�/�.���;�Yt�u�u�u�u����3�_^[�ËD$S3�;�VWt�|$;�w����j^�0SSSSS����������=�t$;�u��ً�8tBOu�;�t��
BF:�tOu�;�u��p���j"Y����3�_^[�U��SV�u3�9]Wu;�u9]u3�_^[]�;�t�};�w�1���j^�0SSSSS�q���������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x��������j"Y���낋L$V3�;�|��~��u��%^á�%��%^�����VVVVV�    ���������^ËD$��t���8��  uP�a���Y�U������   ��3ĉ�$�   �E�SV�u�HW�L$t+Ht$HtHtHtHHtHutj��   �hj�
j�j�j[Q�~WS�:  ����uG�E��t��t��t�d$P���L$P�F����\$@���L$PW�NQPS�D$P�D$$P�:  ��h��  �t$�L<  �>YYt�=H! uV�<  ��Yu�6��;  Y��$�   _^[3�������]�U�����3ŉE�SV3�9�/W��u8SS3�GWhD�h   S�����t�=�/�����xu
��/   9]~"�M�EI8t@;�u�����E+�H;E}@�E��/����  ;���  ����  9] �]�u��@�E �5��3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w��5  ��;�t� ��  �P蔌��;�Yt	� ��  ���E���]�9]��=  W�u��u�uj�u �օ���   �5��SSW�u��u�u�֋�;ˉM���   f�E t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w�5  ��;�tj���  ���P�Ӌ��;�Yt	� ��  �����3�;�tA�u�VW�u��u�u�����t"9]SSuSS��u�u�u�VS�u �l��E�V�����Y�u������E�Y�Y  9]�]�]�u��@�E9] u��@�E �u�:  ���Y�E�u3��!  ;E ��   SS�MQ�uP�u ��:  ��;ÉE�tԋ5��SS�uP�u�u��;ÉE�u3��   ~=���w8��=   w��3  ��;�t����  ���P轊��;�Yt	� ��  �����3�;�t��u�SW��������u�W�u�u��u�u��;ÉE�u3��%�u�E��uPW�u �u��:  ���u������#u�W����Y��u�u�u�u�u�u�����9]�t	�u�����Y�E�;�t9EtP�֊��Y�ƍe�_^[�M�3��l�����U����u�M������u(�M��u$�u �u�u�u�u�u�-����� �}� t�M��ap���U��QQ��3ŉE���/SV3�;�W��u:�E�P3�FVhD�V�����t�5�/�4����xu
jX��/���/����   ;���   ����   9]�]�u��@�E�5��3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w�2  ��;�t� ��  �P�݈��;�Yt	� ��  ���؅�ti�?Pj S������WS�u�uj�u�օ�t�uPS�u����E�S������E�Y�u3�9]u��@�E9]u��@�E�u��7  ���Yu3��G;EtSS�MQ�uP�u��7  ����;�t܉u�u�u�u�u�u���;��tV�ۈ��Y�Ǎe�_^[�M�3��q�����U����u�M�� ����u$�M��u �u�u�u�u�u�������}� t�M��ap���V�t$����  �v�q����v�i����v�a����v�Y����v�Q����v�I����6�B����v �:����v$�2����v(�*����v,�"����v0�����v4�����v�
����v8�����v<�������@�v@�����vD�����vH�߇���vL�ׇ���vP�χ���vT�Ǉ���vX过���v\跇���v`诇���vd觇���vh蟇���vl藇���vp菇���vt臇���vx�����v|�w�����@���   �i������   �^������   �S������   �H������   �=������   �2������   �'������   �������   �������   �������   �������,^�V�t$��t5�;`tP�݆��Y�F;dtP�ˆ��Y�v;5htV蹆��Y^�V�t$��t~�F;ltP蜆��Y�F;ptP芆��Y�F;ttP�x���Y�F;xtP�f���Y�F;|tP�T���Y�F ;�tP�B���Y�v$;5�tV�0���Y^�����U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^��U���S�u�M������]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�o   ��YYt�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�K����� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[��U����u�M��=����E�M����   �A% �  �}� t�M��ap���j �t$����YY�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  �������W�M�E�u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5�N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r;�ur��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC����+�;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5�N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3���A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;�����   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}硠���3�@�   ���e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+���M���Ɂ�   �ً�]���@u�M�U�Y��
�� u�M�_[��U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  �������W�M�E�u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5�N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r;�ur��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC����+�;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5�N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3���A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;�����   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}硸���3�@�   ���e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+���M���Ɂ�   �ً�]���@u�M�U�Y��
�� u�M�_[��U���|��3ŉE��ES3�V3��E��EF3�9]$W�E��}��]��u��]��]��]��]��]��]��]�u軴��SSSSS�    �������3��  �U�U��< t<	t<
t<uB��0�B���/  �$�N��Ȁ�1��wjYJ�݋M$�	���   �	:ujY������+tHHt����  ���jY�E� �  뢃e� jY뙊Ȁ�1���u�v��M$�	���   �	:uj�<+t(<-t$:�t�<C�<  <E~<c�0  <e�(  j�Jj�y����Ȁ�1���R����M$�	���   �	:�T���:��f����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�]���<+t�<-t��`����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*�<	�u��n���j�����J��M��Ȁ�1��wj	��������+t HHt���;���j�����M��jY�@���j�o����u���B:�t�,1<v�J�(�Ȁ�1��v�:�뽃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�[����B:�}��O����M��E�O�? t�E�P�u��E�P�'  �E�3Ƀ�9M�}��E�9M�uE9M�u+E=P  ��  =������  �"��`;��E���  }�ؾx#�E���`9Muf�M�9M���  �E��}���T�����u��q  k�Ƌ�f�; ��]�r��}�����M��u��]��]��S
�M�3��E��EԉE؉E܋¿�  3�#�#�% �  f����<
����  f�����  f������  f���?w3��EȉE���  f��uG�E����u�}� u�}� u	f!M���  3�f;�u!G�C���u9Ku9u�M̉MȉM��  !M��u��E�   �M��U�Ʌ҉U�~U�Lă��M��]��M��U���	�e� �ʋV��
;�r;�s�E�   �}� �^�tf��E��m��M��}� ��]�FF�E��M��}� ����  f��~;�E�   �u-�u؋M��e�������M����ʁ���  f���u؉M��f��M����  f��}B��������E�t�E��M܋]؋U��m�����ًM������N�]؉M�u�9u�tf�M�f�}� �w�Mԁ��� �� � u3�}��u*�e� �}��u�e� f�}���u	f�E� �G�f�E���E���E�f����u�sf�M�f�MċM؉MƋM���M�f�}��f����e� %   � ���e� �Ẽ}� �m����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W�M�_^3�[�6q����V��� �3�x���ė�
���~�-�U���t��3ŉE�S�]VW�u�}�f��U��ʸ �  #ȁ��  f�ɉ]��E���E���E���E���E���E���E���E���E���E���E���E�?�E�   �M�t�C-��C f�ҋu�}�u.��u*��u&f!;f;�����$ �C�C�C0�C 3�@��  f�����   �   �;�f� u��t��   @uh���Qf��t��   �u��u;h���;�u0��u,h���CjP������3���tVVVVV�v������C�*h|��CjP�~�����3���tVVVVV�J������C3��  �ʋ�i�M  �������Ck�M���������ىM�3��"�ۃ�`;�f�U�u�}�f�E��M���  }�x#�ۃ�`�M�;���  �E�T�˃������y  k�M�f�9 ��M�r��}ĥ��Eĥ�MƉE����y
�U�3��Ͼ�  3�#�#��E��E��E�E��� �  f;֍���  f;���  f=����  f=�?w3��E�E�E���  3�f;�u@�E����u9u�u9u�u	f�u���  f;�u$�U�@�B���u9ru92u�u�u�u��  �}�u��}��E�   �U��u�҅��u�~X�T��U��U����U��U��u��6����փe� �4;�r;�s�E�   �}� �}��w�tf��E��m��M��}� �GG�E��M��}� �}���  f��~;�E�   �u-�U��}�u��e������U�������  f���}�U��f��R��  f��}H�����҉U���E�t�E��U��}�u��m�������U�������M��}�U�uσ}� tf�M�f�}� �w�U����� �� � u3�}��u*�e� �}��u�e� f�}���u	f�E� �@�f�E���E���E�f=�sf�U�f�U��U�U�U���U�f�E��f��Ƀe� ��   ��� ���e� �M���k���3��M���f���?��  �H  �u��E��ы�3�#�#�� �  f;Ӎ<�E��E��E�E�����  f;���  f������  f���?w�E���  f;�uG�E����u9E�u9E�u	f�E���  f;�uG�E����u
9E�u9E�t��e� �E��E�   �U��u�҅��u�~R�u؍T��u��U��U��u��6��e� �֋p��;�r;�s�E�   �}� �X�tf� �E��m��M��}� �@@�E��M��}� ����  3�f;�~<�E�   �u.�U��]�u��e����ڋU����ց���  f;��]�U��f;�M����  f;�}B��������E�t�E��U��]�u��m�����ڋU������H�]�U�u�9E�tf�M�f�}� �w�U����� �� � u1�}��u(�}���E�uf�}����E�u	f�E� �G�f�E���E���E�f���rf�ىE�E�Ɂ�   ��� ���M�3��6f�E�f�E��E�E�E���E�f�}���f��Ɂ�   ��� ���M�E�E��E�U��M�f�
t2��M9E'f�" f�}� ��B����$ �B�B0�B ����jY9M~�M�u���j���?  f�E�[�E��}�M��e������E�����K�}�E�uڅ�}2�ށ��   ~(�E�}�M��m�������E������N���}�E�؋E@���Z�]��E���   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B�ҋ�tA�Eȍ0;։U�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K���K�K<5}�M��D�;9u	�0K;]�s�;]��E�sCf� �*؀��ˈX�D �E��M�_^3�[�yh���À;0uK;�s�;ًE�s�f�  f�}� ��@���ʀ��� �P�0�@ �����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u�����   ^t   �3���t��   ��SVW�   t���t   ��t   ��t   ��   �   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#с�   ^[t��   t
;�u �  Ã�@�@�  Ã�SUVW��|$�\$3���tjZ��t����t����t���� t����t��   �ˋ��   #ǽ   �   t =   t=   t;�u��
����   #�t;�u��   ���   f�� t��   �t$(�L$$����#�#��;D$��   ���������D$�l$��|$�\$3���tjZ��t����t����t���� t����t��   �ˋ�#�t$=   t=   t;�u����   ���   #�t��   u��   ���   f�� t��   �T$�=�A ��  �����\$�D$3���yj^f� t��f� t��f� t��f� t��f� t��   �Ƚ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #Ã�@t-�  t��@u��   ���   ���   ��#|$$��#��;�u���   �"���P�D$,�M  Y�\$(�D$(3҄�yjZ�   ��t��f� t��f� t��f� t���   ��t��   ��#�t"��    t�� @  t;�u��   ����#Ã�@t-�  t��@u��   ���   ���   �L$��3���� t   �_^][��������������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ����������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� j
j �t$�  ������U��SVWUj j h���u��%  ]_^[��]ËL$�A   �   t2�D$�H�3���b��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h��d�5    ��3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y��u�Q�R9Qu�   �SQ���SQ���L$�K�C�kUQPXY]Y[� ���U��QQ�EV�u�E��EWV�E��X  ���;�Yu������ 	   �ǋ��J�u�M�Q�u�P���;ǉE�u����t	P����Y�ϋ������@�����D0� ��E��U�_^��jhh�ڊ������u܉u��E���u薞���  �{���� 	   �Ƌ���   3�;�|;�@r!�l����8�R���� 	   WWWWW葰�����ȋ������@��������L1��u&�+����8����� 	   WWWWW�P�����������[P�  Y�}���D0t�u�u�u�u�������E܉U���Ý��� 	   �˝���8�M���M���E������   �E܋U�������u��  Y�U��$������  ��3ŉ�  ��   V3�9�$  �E��u��u�u3���  ;�u'�Z����0�@���VVVVV�    ����������  SW��  �����4��@�����ǊX$������u��]�t��u3��$  ����u&����3��0�՜��VVVVV�    �������0  �@ tjj j ��  �~�������  �N  ��Y�9  ��D��,  ��z���@l3�9H�E���P��4�M�������  3�9M�t����  ����]��E�3�9�$  �E��G  �E��E����=  ��u�3���
���E��ǃx8 t�P4��  ��	  �`8 j��  P�E��P�B�����Yt4�M�+��$  3�@;��V  j�E�SP�
  �������  C�E��jS�E�P��  �������  3�PPj��  Qj�M�QP�u�C�E��l������v  j �E�PV��  P�E�� �4������I  �E��M��9u��E��>  �}� ��   j �E�Pj��  P�E�� ƅ  �4�������  �}���  �E��E��a<t<u�33�f��
��CC�E��u��M�<t<u9�u��0  f;E�Y��  �E��}� tjXP�E��  f;E�Y��  �E��E���$  9E��H����  ���E��T4��D8�k  3ɋ��@��+  �ۋE��M���   9�$  �E��t  ��u��M��e� +M��E�;�$  s'�U��E��A��
u
�E�� @�E��@�E��}�   rы؍E�+�j �E�PS�E�P��4�������  �E�E�;���  �E�+E�;�$  r��  ���E���   9�$  ��  ��u��M��e� +M��E�;�$  s3�U��E��AAf��
u�E�f�  @@�E��E�f�@@�}��  rŋ؍E�+�j �E�PS�E�P��4������$  �E�E�;��  �E�+E�;�$  �p����  9�$  �2  �M��e� +M�j���  ^;�$  s,�U��u��f��
u
f�  �u�u�f�Ɓ}�R  r�3�VVh�  ��  Q���  +��+���P��PVh��  �l���;�tyj �E�P��+�P��5  P�E�� �4�����t	u�;���	���E�;�G�E�+E�;�$  �E��6����0j �M�Q��$  �u��0�����t�E��e� �E��	���E��}� u]�}� t'j^9u�u�җ��� 	   �ڗ���0�6�u�����Y�+�u���D@t�E��8u3��蛗���    裗���  �����E�+E�_[��  3�^�-Z����  ��jh�蟃���E���u�d����  �I���� 	   ����   3�;�|;�@r!�;����8�!���� 	   WWWWW�`������ɋ������@��������L1��t�P�  Y�}���D0t�u�u�u�?������E��辖��� 	   �Ɩ���8�M���E������	   �E�������u��  Y���/h   � x����Y�L$�At�I�A   ��I�A�A�A   �A�a �ËD$���u�<���� 	   3��V3�;�|;�@r����VVVVV� 	   �^�����3�^Ëȃ������@���D��@^ø�á�@��Vj^u�   �;�}�ƣ�@jP�w����YY��0ujV�5�@�hw����YY��0ujX^�3ҹ����0��� ����` |�j�^3ҹ�W�������@����������t;�t��u�1�� B��P|�_3�^��  �=$& t�  �5�0�)Z��Y�V�t$��;�r"��@ w��+�����Q談���N �  Y^Ã� V���^ËD$��}��P胇���D$�H �  YËD$�� P���ËD$��;�r=@ w�`���+�����P�f���YÃ� P���ËL$���D$}�`�����Q�<���YÃ� P���ËD$V3�;�u�;���VVVVV�    �z��������^Ë@^á���3�9�/�����U���SV�u3�;�W�}u;�v�E;�t�3���E;�t�������v�˓��j^SSSSS�0���������R�u�M��'_���E�9X��   f�Ef=� v6;�t;�vWSV�-R�����|���� *   �q���8]�� t�M��ap�_^[��;�t.;�w(�Q���j"^SSSSS�0葥����8]�t��E��`p��u�����E;�t�    8]��0����E��`p��$����MQSWVj�MQS�]�p�l�;�t9]�b����M;�t�������z�H���;��k���;��c���WSV�ZQ�����S���j �t$�t$�t$�t$��������������Q�L$+ȃ����Y�
  Q�L$+ȃ����Y��  U��E�MSVW3��x�E3ۉx�EC���xt�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�&  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP��  �EPSj �u����M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]�U��j �u�u�u�u�u�u�
�����]�U����ESV3ۋ���C��u�t�]tS�%  Y����  �t�Etj�  Y����w  ����   �E��   j��  �EY�   #�tT=   t7=   t;�ub��M�����$��{L�H��M�����{,��$�2��M�����z��$���M�����z��$���$��������   ���   �E��   3��t����W�}�����D��   ��E�PQQ�$�'  �M��]��� �����������}�E���� ��T���]�����Au���3��E�����f�E�����;�}"+��]�t��u���m��]�t�M�   ��m�Hu���t�E����]��E������_tj�   Y�e���u��Et�E tj �x   Y���3���^��[�ËD$��t~���j���� "   ��^���� !   �3��Q��<$�$Y�Q�<$���$Y�U��Q��}��E�M#M��#E�����E�m�E���QQ�L$��t�-L!�\$���t����-L!�$������t
�-X!�$���t	�������؛�� t���$�YY�jh���x��3�9�AtV�E@tH9d!t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%d! �e��U�E�������e��U��x���U�����3ŉE�j�E�Ph  �u�E� �����u����
�E�P����Y�M�3���N����U���4��3ŉE��E�M�E؋ES�EЋ V�E܋EW3�;E�M̉}��}��_  �5���M�QP�օ����t^�}�uX�E�P�u�օ�tK�}�uE�u܃���E�   u�u��k�����YF;�~[�����wS�D6=   w/�������;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P�O��;�Yt	� ��  ���E���}�9}�t؍6PW�u��I����V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u�l���t`�]��[9}ԋl�uWWWWV�u�W�u�Ӌ�;�t<Vj�il��;�YY�E�t+WWVPV�u�W�u��;�u�u��O��Y�}���}��t�MЉ�u�����Y�E��e�_^[�M�3��M����U�����3ŉE��ESV3�9uW�E�N@  �0�p�p�F  ��X���}𥥥�����<�ыH�����Ή}���e� �������ˋ]���׍<;��0�P�Hr;�s�E�   3�9]�8t�r;�r��s3�C�ۉptA�H�H�U�3�;�r;�s3�F���Xt�@�M�H�e� �?�����<��P������Uމ�x�X��4;�U�r;�s�E�   �}� �0t�O3�;�r��s3�B�҉HtC�X�M�E�} �����3��&�H�����P�����������E���  �H�9ptջ �  �Xu0�0�x�E���  ������0�4?�H�����ʅˉp�Ht�f�M�f�H
�M�_^3�[�FK����U���VW�u�M���S���E�u3�;�t�0;�u,�_���WWWWW�    螚�����}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP�|����M������   ���B����t�G�ǀ�-u�M���+u�G�E���I  ���@  ��$�7  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   ���3��u���N��t�˃�0�f��t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �\�]��]ى]��G댨����u�u>��t	�}�   �w	��u,9u�v'������E� "   t�M����E$�����ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^��U��3�9/P�u�u�uuh��P������]ËL$S3�;�VW|[;�@sS������<��@�������@t5�8�t0�=�%u+�tItIuSj��Sj��Sj�� ����3���ȅ��� 	   �Ѕ������_^[ËD$���u蹅���  螅��� 	   ����V3�;�|";�@s�ȃ������@����@u$�y����0�_���VVVVV� 	   螗�������^Ë ^�jh��xq���}����������4��@�E�   3�9^u6j
��w��Y�]�9^uh�  �FP����YY��u�]��F�E������0   9]�t�����������@�D8P����E��8q���3ۋ}j
�v��YËD$�ȃ������@���DP����U�����3ŉE�V3�95�$tN�=t%�u�b  �t%���uf���pV�M�Qj�MQP����ug�=�$u�����xuЉ5�$VVj�E�Pj�EPV��P�l��t%���t�V�U�RP�E�PQ����t�f�E�M�3�^�F������$   ��U���SV�u3�;�t9]t8u�E;�tf�3�^[���u�M��O���E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P������YYt}�E����   ��~%9M| 3�9]��R�uQVj	�p������E�u�M;��   r 8^t8]����   �e����M��ap��Y�������� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p������:����j �t$�t$�t$��������jh���n��3ۉ]�j�9u��Y�]�j_�}�;=�@}W������0�9tD� �@�tP�  Y���t�E��|(��0��� P�X���0�4�2G��Y��0�G��E������	   �E��n���j��s��Y�SV�t$�F�Ȁ�3ۀ�u?f�t9�FW�>+���~,WPV�|���YP�V�����;�u�F��y����F��N ���_�F�f �^��[�V�t$��u	V�3   Y^�V������Yt���^�f�F @tV����P�  YY���^�3�^�jh�m��3��}�}�j��s��Y�}�3��u�;5�@��   ��0��98t^� �@�tVPV�.���YY3�B�U���0���H���t/9UuP�P���Y���t�E��9}u��tP�5���Y���u	E܉}��   F�3��uࡐ0�4�V�-���YY��E������   �}�E�t�E��m���j�^r��Y�j����Y���������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ��U��QQ�E�E�M�]��  ��������f�E��E���U�����U����Dz3��   3�f�E�uc�E�� u9MtU�]��������Au3�@�3���e�E   �t�M�eJ�Et�f�e��;�tf�M ��EQQQ�$�X������%Q���EQQ�$�C����U�����  �����  �E�]�������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��3�PPjPjh   @h�����t%át%���V�5�t���tP�֡p%���t���tP��^�SV�t$W3����;�u�~��WWWWW�    �Ԑ������B�F�t7V�|���V����  V����P�  ����}�����F;�t
P�WC��Y�~�~��_^[�jh0�mj���M��3��u3�;���;�u�~���    WWWWW�R����������F@t�~�E��pj���V�����Y�}�V�/���Y�E��E������   �ՋuV����Y�jhP��i���E���u�}��� 	   ����   3�;�|;�@r�}��� 	   SSSSS��������Ћ����<��@��������L��t�P����Y�]���Dt1�u�~���YP����u���E���]�9]�t�!}���M��}��� 	   �M���E������	   �E��li����u�:���Y�V�t$WV�������YtP����@u	���   u��u�@Dtj�����j�������;�YYtV�����YP����u
�����3�V�<����������@������Y�D0 tW�u|��Y����3�_^�jhp�yh���E���u�>|���  �#|��� 	   ����   3�;�|;�@r!�|���8��{��� 	   WWWWW�:������ɋ������@��������L1��t�P�}���Y�}���D0t�u�����Y�E���{��� 	   �M���E������	   �E��h����u�����Y�V�t$�F��t�t�v�q@���f����3�Y��F�F^����̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[��%��������������hp��K>��Y����̃=�% uK��%��t��%�Q<P�B�Ѓ���%    ��%��tV����i��V蚤������%    ^�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           � � �   $ 6 F X l z � � � � � � � � 	 	 $	 6	 N	 d	 ~	 �	 �	 �	 �	 �	 �	 

 $
 4
 J
 d
 x
 �
 �
 �
 �
 �
 �
  & 4 @ L V b t � � � � � � �   * : L ^ n ~ � � � �         `�        J0R�X�        ����            bad allocation  PolyMass: Vertex Map <-> Polygon Selection plugin v1.2 � 2012 by Keith Young.   v2p.tif res p2v.tif           �?  � � �m �m  n 0 �m  n @n Pn 0n �n �n � �n `n pn 0�   P� .\source\polymass.cpp   Tpolymassexp    h:\maxon\cinema 4d r12\resource\_api\c4d_general.h  %s     h:\maxon\cinema 4d r12\resource\_api\c4d_file.cpp   h:\maxon\cinema 4d r12\resource\_api\c4d_resource.cpp   #   M_EDITOR    T �m             ����MbP?� � 0� � п h:\maxon\cinema 4d r12\resource\_api\c4d_baseobject.cpp h:\maxon\cinema 4d r12\resource\_api\c4d_pmain.cpp  h:\maxon\cinema 4d r12\resource\_api\c4d_basebitmap.cpp �������������h:\maxon\cinema 4d r12\resource\_api\c4d_libs\lib_ngon.cpp  0�h:\maxon\cinema 4d r12\resource\_api\c4d_gv\ge_mtools.cpp   x 	��@	J
�5�5Tv
    e+000      �~PA   ���GAIsProcessorFeaturePresent   KERNEL32    CorExitProcess  mscoree.dll .mixcrt EncodePointer   KERNEL32.DLL    DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    X'�'runtime error   
  TLOSS error
   SING error
    DOMAIN error
      R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:                      �?5�h!���>@�������             ��      �@      �            	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ =    Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        ������x�l�`�T�L�@�4�
�x�\�H�(��,�$�� ������ ���������������������������������������������������������������x�l�d�X�@�4� � ���������\�@����������������h�`�T�D�(��������d�H�$� �������
�InitializeCriticalSectionAndSpinCount   kernel32.dll    ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx          GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL                                                                                                                                                                                                                                                                                        ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun 1#QNAN  1#INF   1#IND   1#SNAN  _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   modf    fabs    floor   ceil    tan cos sin sqrt    atan2   atan    acos    asin    tanh    cosh    sinh    log10   log pow exp SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    CONOUT$     ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           ��              h�t���           ����    @   X�         ����    @   ��           ����               ����t���    8       ����    @   ��            P            $ 8 ��t���    P       ����    @                 ��           x �     �        ����    @   h             ��            � �     �        ����    @   �             ��            �     �       ����    @   �             D           T\            ����    @   D            0�           ��    0        ����    @   �            P�           ���     P       ����    @   �            t            08    t        ����    @                �h           x�    �        ����    @   h    p7 �p ��                     ����    ����    ����>O    ����    ����    ����    �    ����    ����    ����        ����    ����    ����    /    ����    ����    ����    �"    ����    ����    ����    �%    ����    ����    ����    �(    ����    ����    ����    D*����    P*����    ����    ����Y/]/    ����    ����    ����    �;    ����    ����    ����    z=    ����    ����    ����yQ�Q    ����    ����    ����    �T    ����    ����    ����    �X    ����    ����    ����    \    ����    ����    ����9iMi    ����    ����    �����i�i    ����    ����    ����    }k    ����    ����    ����il�l    ����    ����    ����    �m    ����    ����    ����    o    ����    ����    ����    1�    ����    ����    ����    /�    ����    ����    ����4�P�    ����    ����    ����    �    ����    ����    ����    ��    ����    ����    ����    F�        �����    ����    ����     �    ����    ����    ����    ��    ����    ����    ����    F��         �  �                     � � �   $ 6 F X l z � � � � � � � � 	 	 $	 6	 N	 d	 ~	 �	 �	 �	 �	 �	 �	 

 $
 4
 J
 d
 x
 �
 �
 �
 �
 �
 �
  & 4 @ L V b t � � � � � � �   * : L ^ n ~ � � � �     FGetCurrentThreadId  GetCommandLineA HeapFree  �GetVersionExA HeapAlloc �GetProcessHeap  qGetLastError  �GetProcAddress  GetModuleHandleA  � ExitProcess eTlsGetValue cTlsAlloc  fTlsSetValue dTlsFree ,InterlockedIncrement  (SetLastError  (InterlockedDecrement  VSleep $SetHandleCount  �GetStdHandle  fGetFileType �GetStartupInfoA � DeleteCriticalSection }GetModuleFileNameA  � FreeEnvironmentStringsA UGetEnvironmentStrings � FreeEnvironmentStringsW �WideCharToMultiByte WGetEnvironmentStringsW  HeapDestroy HeapCreate  �VirtualFree �QueryPerformanceCounter �GetTickCount  CGetCurrentProcessId �GetSystemTimeAsFileTime ^TerminateProcess  BGetCurrentProcess nUnhandledExceptionFilter  JSetUnhandledExceptionFilter 9IsDebuggerPresent HeapSize  QLeaveCriticalSection  � EnterCriticalSection  �VirtualAlloc  HeapReAlloc �WriteFile GetCPInfo � GetACP  �GetOEMCP  ?IsValidCodePage RLoadLibraryA  #InitializeCriticalSection �RtlUnwind uMultiByteToWideChar tGetLocaleInfoA  DLCMapStringA  ELCMapStringW  �GetStringTypeA  �GetStringTypeW  SetFilePointer  "GetConsoleCP  3GetConsoleMode  �RaiseException  7SetStdHandle  �WriteConsoleA 5GetConsoleOutputCP  �WriteConsoleW S CreateFileA 4 CloseHandle � FlushFileBuffers  KERNEL32.dll                    ���O    "              `�  /   PolyMass.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         `�`���    .?AVNodeData@@  ��    .?AVBaseData@@  ��    .?AVTagData@@   ��    .?AVPolyMass@@  `�`�`�`�`�`�`�`�`�`�`�`���    .?AVGeSortAndSearch@@   ��    .?AVNeighbor@@  ��    .?AVDisjointNgonMesh@@  `�`�`�`�`�`�`�`�`���    .?AVGeToolNode2D@@  ��    .?AVGeToolDynArray@@    ��    .?AVGeToolDynArraySort@@    ��    .?AVGeToolList2D@@  `�            u�  s�  `���    .?AVtype_info@@ N�@���D    sqrt    �g�g�g�g�g�g�g�g�g�g`�            �%��������    �����
                                                                   �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �             x   
                                                                                                                                                                                                                                                                                        ��   t�	   H�
   ��   ��   T�   0�   �   ��   ��   l�   4�   �   ��   ��    P�!   X�"   ��x   ��y   ��z   ���   ���   p�                                 	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                               ���5�h!����?      �?                                                                                                                                                                                                                                                                                                                                          abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     p�  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    L�����C                                                                                              �            �            �            �            �                              `        H���P���   �p        p�`�H�J�x�t�p�l�h�d�`�X�P�H�<�0�(�������� ������������������������������������|�p�\�P�	         �.   \�/�/�/�/�/�/�/�/�/`   .         ���5      @   �  �   ����              �            �0    �0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                `�   \�   X�   P�   H�   @�!   8�   0�   (�    �   �   �   �   �    �   ��   ��   ��   ��   ��   ��   ��   ��   ��"   ��#   ��$   ��%   ��&   ���&         �D        � 0     �p     ����    PST                                                             PDT                                                             x!�!����        ����                 �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                 �      ���������              �����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l  ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �                 0  �              	  H   XP V   �      <assembly xmlns="urn:schemas-microsoft-com:asm.v1" manifestVersion="1.0">
</assembly>PAPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDING   �   00P0^011�1�1�12i2�2�2�2�2�2313x3�3�3�3�34=4�4�4$5t5�5$6>6]6�6�6�6�667a7�7�7�7�9�9C:]::�:�:�:;;);L;y;�;�;�;�;<$<5<T<q<�<�<�<�<$=A=d=�=�=�=>4>d>�>�>�>?$?D?d?�?�?�?�?�?      �   0!010D0d0�0�0�011$1d1�1�1�1�122!242T2t2�2�2�2�23D3d3�3�3�3�3�34?4a4t4�4�4
545T5t5�5�5�5�5646T6t6�6�67T7�7�78T8�8�8�89!949d9�9�9�9�9�9:$:D:d:�:�:;(;E;h;�;�;�;<2<F<V<�<�<�<�<�<=4=T=t=�=�=�=�=>=>R>t>�>�>�>�>?$?>?R?b?�?�?�?�?�? 0    0!0O0t0�0�0�0�011D1\1�1�1�1�1�12=2k2~2�2�233T3t3�3�3�34$4D4d4�4�4�4�4�45D5d5�5�5�5�56$6D6d6�6�6�6�6�6�6$7A7Q7t7�7�7�7�7�7�788,8Q8t8�89D9t9�9�9�9�9�9:%:3:T:e:s:�:�:�:�:;!;1;T;l;�;�;�;�;�; <<<0<T<l<�<�<�<�<�<�<!=1=D=d=�=�=�=�=>>'>D>t>�>�>�>??4?a?t?�?�?�?�?   @    040T0q0�0�0�0�0�01$1D1d1�1�1�1�1�12D2^2u2g3�3�3�3�3�3�3�4�4�4�45D5d5�5�5�5�56$6D6a6t6�6�6�6�6717D7_7m7{7�7�7�7�7�7 8!8D8d8�8�8�8�8�8�8�89/9=9K9Z9l9�9�9�9�9:4:T:t:�:�:�: ;;-;W;i;�;�;�;�;�;<4<T<t<�<�<�<�<�<�<=4=N=b=q=�=�=�=�=�=>,>=>K>b>w>�>�>�>�>�>??&?q?�?�?�?�?�? P    0$0D0d0�0�0�0�01$1D1d1�1�1�1�12$2D2d2�2�2�2�23@3d3�3�3�3�34$4D4d4�4�4�4�45$5D5d5�5�5�5�56$6D6d6�6�6�6�6�6717D7a7q7�7�7�7�7�7
88D8d8�8�8�89"9:4:N:^:o:�:�:;4;Z;h;w;�;�;�;7<k<�<�<�<===4=A=N=f=y=�=�=�=�=�=�=>">8>T>e>x>�>�>�>�>�>�>??(?F?d?v?�?�?�?�?�?�?   `    000F0b0s0�0�0�0�0�0�011/181V1t1�1�1�1�1�1�122@2V2r2�2�2�2�2�2�23D3R3_3w3�3�3�3�3�3�34424H4d4v4�4�4�4�4�455&5/5M5n5�5�5�5�5�5�56,6W6�6�6�627:7D7V7`7{7�7�7�7�7�7/8M8v8�8�8%979H9Q9d9�9�9�9:(:::L:r:�:�:�:t;�;�;<D<R<q<�<�<�<�<=!=4=T=t=�=�>�>?�?   p  �   000%0,030:0A0H0O0V0]0d0k0r0y0�02A2l2�2�2�2C3U3�3�394U4�4�495\5x5�5�5�5�56}6�67l7�7�7848T8t8�8�8�8�8949T9q9D:r:�:�:;R;�;�;%<U<e<�<�<A=}=�=>E>�>�>�>5?u?�?�? �  �   E0�0�0�0%1b1�1�12e2�2�2%3h3�3�3�3�3�3E4�4�45E5�5�5"6q6�6�6�6�6 7%7M7t7�7�7�7%8I8�8�89)9R9�9�9�9:H:�:�:�:;�;�;�;�;<$<D<a<�<�<�<�<=4=T=q=�=�=�=>�>�>!?A?a?�?�? �  �   $0t0�0�0�0141T1t1�1�1�1�1$2D2t2�2�2�2343a3�3�3�3414T4�4�4�4515Q5q5�5�5�5�5616Q6q6�6�6�6�6717Q7t7�7�7�7848a8�8�8�8�89A9d9�9�9�9:^:�:�:�:;$;D;t;�;�;�;<!<D<t<�<�<�<=D=d=�=�=�=�=>$>A>q>�>�>?d?�?�?�?�?   �  �   0D0q0�0�0�0111Q1q1�1�12$2T2�2�2�23D3�3�3�3!4A4a4�4�4�455545]5�5�5
646T6z6�6�677�778q8�8�8�8�89=9s9�9�9:!:D:d:�:�:`;�;�;�;<4<i<�<�<�<�<=2=S=t=�=�=�=>1>T>t>�>�>?4?a?�?�?�?   �  �   0040�0�0�0141T1�1�1�1�1A2^2�2�2�2�23;3L3l3�3�3�3�34.4B44�4�4�45;5S5q5�5�5�5�5�6�6�6�677?7d7�7�9�<�<�<=F=V=�=�=�=�?�?�?�?�?   �  �    0{0�0�0�0!1(1/1�1�1�1�1�1$2D2t2�2�2�233D3d3�3B4H4v4�4�4�4�4�4�4(5;5U5l5p5t5x5|5�5�5�5�5�56A6�6�6�6�6717D7t7�7�7�78$8D8t8�8�8�8949T9t9�9�9:(:7:t:�:�:�:;1;T;t;�;�;�;<1<�<�<�<4=Q=d=8?J?]?�? �  `   N0f0�1!242d2�2�2�2�23333T3t3�3�3�34%444a4�4�4�4�4�4$5T586l6�6�6;788&8�8�8�8B9�9�9   �      ?4�=>->e>�>�>5?u?�?�?   �  p   "0U0�0�01E1�1�1222b2�2�2�253u3�34U4�4�45e5�5%68+8�:8;<;@;D;H;+<9<X<f<�< =%=-=�=�= >.>g>u>|?�?�?�?     �    0.0C0Q0W1h1:5�5�5,7`7�7�7�7858H8o8�89�9�9�9�9�9 ::
:::::#:':-:1:7:;:A:E:Z:k:�:�:�:�:;;,;1;7;=;i;n;x;�;�;�;�;<"<=<n<�<�<�<"=�=�=�=>7>b>g>|>�>�>'?1?R?�?�?�?�?  �   =0C0T0r0�0J11�1�1�1�1�1�1�12!2(2,2024282<2@2D2�2�2�2�2�233,33383<3@3a3�3�3�3�3�3�3�3�3�3�3*4044484<4�4�4"5-5?526=6j6r6�6�669�9�9#?�?   d  z1�1�1�1�122$2D2I283M3S3\3c3�3�324:4F4N4b4m4r4�4�4�4�4�4�4�4�4�4555Y5^5i5n5�566N6g6�6�6�6�6�6�6�6�6
777'7<7B7V7]7w7�7�7�7�7�7�7�7�7�7�7�7�7�7 88%8.8;8\8f8�8�8�8�8�899>9�9�9�9::^:q:w:�:�:�:�:�:�:�:�:�:�:�:�:�:;
;;;;$;,;5;A;F;K;Q;U;[;`;f;n;z;�;�;�;�;�;�;�;�;�;�;�;<<0<_<h<t<�<�<�<�<�<==3=T=Z=�=�=�=+>5>]>v>�>�>�>K?Q?s?�?�?�?�?   0   	00^0i0q0�0�0:2M2U2[2`2h2�2�2�2�233&3-3d3�3�3�34 4%4D4I4�4�4�45	555)525;5M5V5b5k5r5|5�5�5�5!6'6@6F6	7&77c8k8�8�8�8909=9I9Q9Y9e9�9�9p:v:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;
;;!;&;6;;;A;G;];d;m;�;�;�;<<#<M<Y<_<�<�<�<�<�<�<�<�<�=�=�=�=�=�=�=�=�=�=�=>   @ �   D0R0X0r0w0�0�0�0�0�0�0�0�0�0�0�0111$1,121<1C1W1^1d1r1y1~1�1�1�1�1�1�1�1?2�5�56<6v6�6�8�8�8�8�899>9G9N9W9�9�9�9�9::7:I:n:�:�:�:�:;;F;T;w;<</<�=0>�>L? P �   011-151E1V1_12�2�2�2^4o4�4�4�4�4�4�455(5A5K5^5�5�5�5�5o6�6�667U7�7�7�7�788&8=8V8r8{8�8�8�8�8�8�8�89�9
:T:�:�:";�;�;�;�;<)<�<�<�<�<�<=�=�=�>�>�?   ` �   j0�0�0�0�0�0�0�0�0#1A1H1L1P1T1X1\1`1d1�1�1�1�1�1&212L2S2X2\2`2�2�2�2�2�2�2�2�2�2�2 3J3P3T3X3\36�8�8�8�8�89n9�9�9�9�9�9�9�9::Y:^:�:�:�:�:�:�:/;8;>;�;�;�;�;�;(<.<7<><I<U<�<�<==b=h=t=�=�=4>�>�>�>�> ?C?w?}?�?�? p h   ]0i0u1�2�2�3a4y4�4�45)5A5�7�8�9�9�9�;==== =$=(=,=2=J=a=g=w=|=�=�=�=�=�=�=�=�=
>>>*>�>�>�> � l   /060<0�0G1}1�1�1�1�1�1�1�1%2�2k3�34�4a5k5�5�5�5�5�5�5�5y6�6�89919C9U9g9y9�9�9�;�<�<e=G>�>�>�?�?�? � T   >0U0�0�1�1�2�3"4(4�4�4�4�5�5�5R6"999N<R<V<Z<^<b<f<j<n<r<v<z<�<[=s=�=�=>2>   � 0   �7t:�:�:];w;�;�;�;<%<c<�<J=�=c>�>X?~?�? � �   �0�1P2w2�2�2�2`3�3�3;4�4�4�4�4�455&545;5J5V5c5�5�5�5�5�5�56!6*6M6w6�6�6�7�7�:�;<#<9<A<�<�=�=�=
>>%>U>�>�>�> ??�?�? � �   y0p4�4�4�4�4�4<5M5�5�5�5	636A6M6[6c6p6�6�6�6�6�6�6�6�6�6�7858V8b8�8�8�8�8x9�9�9�9:�;�;�;�;�;
<�<=:=b=�=�=><>F>^>�>�>�>   �    P0a0r0z0�0�0�0�0 � p   $1014181<1@1L1P1�1�1�1�1�1�1�1�1 22222222 2$2(2,20233034383<3@34484x4|4�4�4�4�4�4�4�4�4�4h5l5   � �   �1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,2024282<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3L?P?d?h?l?t?�?�?�?�?�?�?�?�?�?�?�?     �   00 0$0(0,00080P0`0d0t0x0�0�0�0�0�0�0�0�0�0�01111,1<1@1P1T1\1t1�1�1�1�1�1�1�1�1�1�1�1�1222,20282P2`2d2t2x2�2�2�2�2�2383X3x3�3�3�3�3�3 4 4<4@4`4�4�4�4�4�4�4 55 5@5`5�5�5�5�5�5 6 6,6H6h6�6  0   000 080P0h0l0p0t0x0|0�0�0�0�0�0�0�0�0�0�0�0�0�0 11111101P1t1�1�1�1�1�1�1�1�1�1�1�1�1�1 2244$4,444<4D4L4T4\4d4l4t4|4�4�4�4�4�4�4�4�4�4�:�;�;<<(<8<\<h<l<p<t<x<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$=(=,=0=4=8=<=@=D=H=X=`=d=h=l=p=t=x=|=�=�=�=�=�=   H   d0l0t0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01111$1,141<1D1�1�1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              