MZ�       ��  �       @                                      � �	�!�L�!This program cannot be run in DOS mode.
$       �CZʍ"4��"4��"4���"4�|����"4�|����"4�|����"4��"5��"4�qU���"4������"4�/����"4�/����"4�/����"4�Rich�"4�                        PE  L `�
R        � !  J  �      ^�     `                         p                             �� K   �� (                            @ �   Pa 8                            � @            `                           .text   %I     J                   `.rdata  �   `  �   N             @  @.data   �1         �             @  �.reloc  �-   @  .   �             @  B                                                                                                                                                                                                                                                                                                                                                                        V����\  ��aW��N8�N@�NH�NP�NX�N`�Nh�Np�Nx���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ��   ��  ��  ��  ��   ��bf֎(  fֆ@  f֎X  f֎p  f֎0  f֎H  fֆ`  f֎x  f֎8  f֎P  f֎h  fֆ�  f֎�  fֆ�  f֎�  f֎�  f֎�  f֎�  fֆ�  f֎�  f֎�  f֎�  f֎�  fֆ�  f֎�  fֆ   f֎  f֎0  f֎�  f֎  fֆ   f֎8  f֎�  f֎  f֎(  fֆ@  �F    �F    �F     �F(    �F,    �F0    ǆd      ǆh      ǆl      ǆp      ǆt      ǆx      ��^���������V����a�rI  ��^�JZ  ����������U��VW�u�}�u��W��  ����u_3�^]� �M�F ǆd      ǆt      f�F �j �@h�  ���   ��j �΃�uWj W�  ������t��W�@H�v��$  ���~ f�FP�~@��f�FX�~@_f�F`�F�   ^]� jW�  �������H���_�F �   ^]� ����������U��V���eH  �u���u��  ^]� ���U���dS�]W����u
_3�[��]� ����t  ��t_�   [��]� S����  ������tɀ V��   � ��   � ��   ��P  ���   �O0�E�P� M  �O0���&M  ��P  �v�F0�^ �I�N(���l��d����Y��Y��Y��Y��X6�X^j �XNh �X��FH�Y��X��F8�Y��X��FP�Y��X��F@�Y��X��FX�Y�f�wPf�_X�G�X�f�O`��  ���G ^_�   [��]� hN� S���  ���E���tP����u  ����t@3�9w$t)3ۋG�Mj �4j(��u  ����tF��;w$u܋]����u  ����u^_3�[��]� �u���u�u�u�S�J$  ^_[��]� �U��V�u��u3�^]� ���s  ��u�W���   ���   �ЉE��tcjP����a  ��M���   ���   �Ћ�3���t;�V���   �M���   �Ћ�Ћ��   h$  �@���Ѕ�u*F;�u�3���E���   P���   �у���_^]� �   @����������U����0�@V�@ W�}$�����=mric��  hv'  ��  ����RP�B8j���Ѐ~ ��  �}W�u��f�F  �F ��  �E�\F8���   �\N@�E��E�\F@�M��E����   �\F8�E��^��o �E��r �E��E��St �]�f(��YE�f(��Ye�f(��YM��YU��\�f(��Y]��YM��\��\�� cfTcf/�v?W�f/�vf/�vf/�wf/�v$f/�vf/�v���F��  _�   ^��]�  ���   �\F8���   �\N@�E��^��M���n �E���q �E��E��ys �]�f(��YE�f(��Ye�f(��YM��YU��\�f(��Y]��YM��\��\�� cfTcf/�v?W�f/�vf/�vf/�wf/�v$f/�vf/�v���F�"  _�   ^��]�  ���   �\F8���   �\N@�E��^��M���m �E���p �E��E��r �]�f(��YE�f(��Ye�f(��YM��YU��\�f(��Y]��YM��\��\�� cfTcf/�v?W�f/�vf/�vf/�wf/�v$f/�vf/�v���F�H  _�   ^��]�  ;�t  t�F�~ ��   �E�P�E$P�E�P�EP��辙  �E�+E�}$+}@�E썆d  PG���  ��詜  ��d  ��u
_3�^��]�  ��M�@j ���   h�  �Ћ�d  j Pj�v �u�u�W�!�  ����t��E�F ��t  �,E��P�,EǆP  ����P��  ���g  _�   ^��]�  ����������U��V�uWV�u�����  �j �@h�  �@0���Сj�@h�  �@4�����G _^]� �������U��E���  S�٨��
  ���
  V�uV�  ������u^[��]� �{ u
f�C  �C WV�u����  �}WV���  ��bW������j/P��p�����x����E���X�����`�����h����E��E��M���0�����8�����@���较  ���{ ��  ��`  �� �  H��   H�  ��b��bfօx���f�E�fօX���fօh�����bf֍p���f֍`�����bf�E�f�E���bf�M�fօ0���fօ8���f֍@����  ��b��b��b��bfօX���fօh�����bf֕p���f֍x���f�M�f֝`���f�M�f�M�f�U�fօ0���f֝8���fօ@����  ��b��b��bfօx���f�E���bfօ`���f�E���bf֕p���f֍X���f֍h���f�M�f�M�f֕0���fօ8���fօ@����   �{ t/�~����fօp����~� ���fօx����~�(���f�E��e�{ t2�~����fօX����~� ���fօ`����~�(���fօh����-�{ t'�~����f�E��~� ���f�E��~�(���f�E���M��E�   �E�   �@dQ���   h�  W�С�M؋��   Q� �Сj �@d��p����@QW�С�s8�Hd���   P�A$VW�Сj �@d��X����@QW�С�Hd���   P�A$VW�С��@�@dj �@�M�QW�С�Hd���   P�A$VW�С�M��E�   �E�   �@dQ���   h�  W�С�M؋��   Q� �Ѓ�(�{ u	�C�   ��P  ���   �������@HQ�K0�@,�Ћ��   ��p����@d�}�@p��p���Q�s0W�Сj�@dW�@`�Сj �@d������@QW�ЋK0�� �B  ��P  j �Ij�ȡQ�@dW���   �Сj �@dW�@`�Ѓ��{ ��  ��`  W�f(�f(�f(���P�����H����u��E��E��E��� ��   HtxH�O  ��b��E��E��M��@dj �@�M�QW����b���   �ch�kp�sx�Y��M����   �Y��M����   �   ��b��E��M��Eȋ@dj �@�M�QW���ch�kp�sx�C��b��M��E��E��@dj �@�M�QW�����   ���   ���   ��b���   �Y��M����   �Y��M����   �Y��Y��Y��Yȃ���P�����H����u��M��[P�SX�K`(��\��X܍E�P�������E�(��\��X�P���]��E�(��\��X��U��E��M��;@  ���E�P�� ���P���'@  �V�IdP�A$W���[P�SX�K`f(��\E��X]����E�P�E�f(��\E��XU��� ���P���E�f(��\E��XM��]��U��E��M��?  ���E�P������P���?  �V�IdP�A$W����  �X[P�SX���X�  ��   �XK`f(��\�P����X�P����E�P�� ����E�f(��\�H����X�H���P���]��E�f(��\E��XM��U��E��M���>  ���E�P������P����>  �V�IdP�A$W����  �X[P�SX�X�  ��   �XK`f(��\E��X]����E�P�E�f(��\E��XU��� ���P���E�f(��\E��XM��]��U��E��M��L>  ���E�P������P���8>  �V�IdP�A$W�Ѓ���  �XCP�E�P������P�E��CX�X�  ���E���   �XC`�E���=  ��������@dQ�@$�K8QW�С�M��E�   �E�   �@dQ���   h�  W�С�M؋��   Q� �Сj �@d��0����@QW�Ѓ�(�{ ��   ���   V�� ���P���O=  �P�Id������P�A$W�Ѓ�������8  �P�Idj �ApW�Сj�@dW�@`�Сj �@d������@QW�Сj �@dj���   VW�Сj �@dW�@`�Ѓ�8�Ffn�X  �����M��E�fn�\  ���Q�E�W��E��@d�������@$QW�Ѓ���M��E�   �E�   �@dQ���   h�  W�С�M؋��   Q� �Ѓ�_^�   [��]� 3�[��]� �����������U��S�ًMj � �  �8�  u&��M�@j ���   h�  �Ѓ�t3�[]� �u���u�u�u�u�u���  []� ����U��}S�]VW�}��uqW�  WS���	  �j �@h�  ���   ���Ѓ�u@�~ u>�W�@H�v��$  ���~ f�FP�~@f�FX�~@��f�F`�F��F �u���uSW��  _^[]� �����V��P  ;�T  u�F:Fu�F:Fu�F:Ftj h �F��v  ���F �F�F�F�F�F�F��P  ��T  ^��������������U����  �} S��u.����   ���   �ЉE��u	2�[��]� �MjP�`P  ����   ���   �ЉC ��tҡ�M���   ���   �ЋЉU̅�t��h`b�H�R��h�  P���   �Ѓ��C��t�W3��} �C$    �}�tW�f�KPf�KXf�K`V3��u����M���   V���   �Ћ�Ћ��   h$  �@���Ѕ��P  ��M���   W����   Vf�E�f�E�f�E��ЋЉS�R���   �K ���   �ЋC$�K�@�C�ыK�:�  �K$�I�K�D��C$�@�C�L��Q�@\�@X�ЋK$���I�K�D��C$�K�@�L���  �K$j �I�Kh�  �D���s�@H��p  �ЋK$���I�K�D��C$�@�C�L����N  �h`b�@�����   h�  Q�ЋK$���I�K�D��C$�@�C�|� ��  �K�E�P�E�P3�h���V3��u�E�  ���.�  �} �=  ����   G�}�}�;}���   ������E��C$�K�EЍ@�E�D�E��� �X �E��@�XE��E��@�D��XEĉ|��C$G�@�C�EċT�U��D��E��~f�D0��~Bf�D0��~Bf�D0�;}��t����u�}�K�E�P�E�Ph���W�h�  ���Q�  ���-����}��} ��  ���<����@HQ�K�@,�Ћ��C$�   ��������������@�CfnD������@H�Yȋ@,������Q�K�M�������Y��M�������Y��M����m��e��uċ�   ��\������t����]��U��Y��Y��M��Y��X��E��Y��Y͋}��X���|����Y��X]��X��E��Y��X[P�X��E��Y��[P�XU��X��E��Y��XSX�X��SX�XM��XK`�K`�C$�@�C|��}��   ����   G�}�}�;}�k������E���$    �C$�E�@�C�v �D��|��C$G�@�C�T�U��D��E��~f�D0��~Bf�D0��~Bf�D0�;}�~��u�}�K�E�P�E�Ph���W�_�  ���H�  ���a����}��C$�u�F�u�;u��j����} t\fn����W�f.����D{8��b�^��CP�Y��CP�CX�Y��CX�C`�Y��C`��K`�KX�KP��M���   Q���   �Ѓ��{$ u^_2�[��]� �C��������K�R�@H�@,��W���(  ��   �fփ�   fփ�   fփ�   f�C8^fփ�   fփ�   fփ�   f�C@_fփ�   fփ�   fփ�   f�CHf�C  �C ǃP  ����f�C  �C �C ǃd      �C0    �C �[��]� ������U����V���   �񋀈   �u��ЉE��u	2�^��]� �MSWjP�I  ��M􋀈   3ۋ��   �б3��E�M�����   3����    ��M􋀈   W���   �Ћh$  ���   �ȋR�E��҅�t7�E�;X$}i�H�E��;u]��q�@\�@X�ЋM����I9D1u>C��G;}�u��M��u�;^$_[u+��t'��M􋀈   Q���   �Ѓ��^��]� 2��ˋ���,  �u��j �u����^��]� ��������U����ESV��E��E3�ǆp      �E�� �E�9^$tlW3���d  j j j j�E�P�E�P�F�48�N�  �E���t7�U��M�+M+U�����;M�}��p  �F�M��F0�E��@��P  C��;^$u�_^[��]� ��������������U����   �@S���   V�uWj ��h�  ����H���%  �$�x1 �������*-  ���  ��K���   �@0�Ћ�����   ����   �΋R0�ҋЅ�t(���$    �d$ ��򋁈   �ʋ@0�ЋЅ�u��M��@HQ�@,���Ћ��   ��K���   �@0�ЋЅ�uF��@����,  ���r�M��\  �P�Ih�E�P�A�Ѓ����P�u��h�  �>  �Ѕ�t5��AH�M��@,Q���Ћ��#��u�@H�s��$  �Ѓ������(  ���  W����   �f�R��@���f�BPf�B�4,  �����  �   ���_^[��]� �0 )1 0 �0 �0 �0 1 ������������U���   ��bSVW�}�E�P�E�P�E�P�ٍE�P����H  舁  �u�+u�W�+u���p���u�P�E�P��X���P����X�����`�����h����E��E��E���p�����x����E�脁  �W�@h�@�Ѓ����  �E��M�+E�+M�;�~fn��fn������@h�KP�@8Q�M�WQ�E����u�~ f�E��~@f�E��~@�W�@d�E��@X�Ћȃ���u�W�@d�@�Ѓ��ȡQ�@@�@,�Ћ�c�QQ���   ���$h�  �����]���c�@�����   �$h�  �����]��E��^Eȋ}�YE�fn�����Y��^E��fn�����^E��Y�H  �sPV�M���H  �W�@hQ�@,����H  �~ f�C8�~@f�C@�~@f�CH���  ���  W��Y��Y����  f(��Y��  �X����  �Y��Y��X����  �Y��X����  �Y��X����  �Y��X����  �Y�f�[hf�Sp�X�f�Kx���  ���  ���  �Y��Y��Y�(��X����  �Y��Y��  �X����  �Y��X����  �Y��X����  �Y��X����  �Y�f֛�   f֓�   �X�f֋�   ���  ���  �Y��Y��X�(��Y��  �X����  ���  ���  �Y��Y��Y͍M��X����  �Y��Y��  Q�X����  �Y�f֛�   f֓�   �M��X�WQ�X�f֋�   �Ch�X��E��Cp�XF�E��Cx�XF�E�@h�@,���~ fփ�   �~@fփ�   �~@fփ�   ���   �X��M�Q�M��E����   �XFWQ�E����   �XF�E�@h�@,���~ fփ�   �~@fփ�   �~@fփ�   ���   �X��M�QW�E����   �XF�M��E����   �XF�E�@h�@,Q���~ fփ�   �~@��0fփ�   �~@_^fփ�   [��]� ����������U�������   V���   ���Љ�x  ��u	2�^��]� �MSW��>  P���  �M�E�P�E�P�E�P�E�P�'|  �}��]�+}�+]�GC�$  ��h  ��tw���x  ���   ���   �Ѕ�t&��h  j �uj��x  �uSW�  ����t4�} t9��~  ��l  ��tj �u��j�v �uSW�l  ����u_[2�^��]� _[�^��]� �������������V��h  P�~  ����   ��x  P���   �Ѓ�^��̍�l  P�T~  Y���U��SW�}�م���   V�W�@@�@�Ѓ����   �j �@HW���   ���Ѓ���t2�j �@HW���   �Ћ������   �΋@4��P���   �V�@H���   �Ѓ���t�V�@H���   �Ѓ�����x  ���   V���   �С�ϋ��   �@4��P���$�����ϋ��   �@(�Ћ�������^_[]� �U��SV�u�م��   W�V�@H�����   �Ѓ���t�V�@H���   �Ѓ����W���   ��x  ���   �С�΋��   �@4��P��������΋��   �@(�Ћ���u�_^[]� ���������U���4  S�ـ{ tǃ`      �"�{ tǃ`     ��{ t
ǃ`     �~CPf�E��~CX�Mf�E��~C`f�E��~CPfփ�   �~CXfփ   �~C`fփ  W�fփ  fփ  �C�C fփ   �j �@h�  ���   ��jP�u���u�>���������u�ˈC�H!  3�[��]� VW��������3  ��M�@3����   Whxvpi�E� ǅH���    ǅ\��������}��ЋM��X  �W�@hyvpi���   �Ћufn����j�����D$fn�X  �����\  �$h �  �t�  ������P��8���P��0���P��蘽  ����  �j �@haqpi���   ����������0�����8����ȃ�W�f.Љ�l������Dzf.ȟ��Dz;��  �}� tw��h  P�z  ����   ��x  P���   �С�M�@�����   j h�  ��j P�u���u�����������(  ��8�����0����E� fn�X  ���ǃp      �X¿�� �}3��,�fn�\  �����X  �X���p�����x  �,���\  ��h�������   ���   �Ѕ���   ��    ���x  ���   V���   ��j j j j��h���Q��p���Q��h  P�E�z  ��t2��h�����p���+�X  +�\  �����;�}��p  �E���C(���x  ���   F���   ��;��i����}3��E�����9s$tv3���    ��l  j j j j��h���P��p���P�C�4�z  ��t:��h�����p���+�X  +�\  �����;U}��p  �C�U��C(�u�F��;s$u���p  ���3  ��H���9K(u��\���9Hu�}�9�l����$  ��^  ��������@Q�@�Сj �@j��@������h�bQ�Ћ�p  �H�Q�@�������@(Q�Ћ���I�������IP�ы�A�������@QV�С�������@Q�@�С�K(���   ��,�@x��hw'  ���h�  ����I������IP�ы�A������@QV�С���@������@<�Ћj��Qj�WP������BL��hx'  ��  ����I�� ����IP�ы�A�� ����@Q�����Q�С���@�� ����@<�Ћj��Qj�VP�BL�� ����С�������@Q�@�С�������@Q�@�� ���Q�С���@�������@<�Ћj��Qj�������QP�BL�������С�� ����@Q�@�С�� ����@Q�@������Q�С���@�@<�� ����Ћj��Qj�������QP�BL�� ����Ѝ� ���P��\  ��� ����@Q�@�С�������@Q�@�С�� ����@Q�@�С������@Q�@�С�������@Q�@�С�������@Q�@�Ћ�p  �K(�C�B��\����E�����H����K,����^  �r�4@�C���u��L�Q�@\�@,�Ѓ����2  �~CP�Cfփ�   �~CXfփ   �~C`fփ  �T3ɉM����  ��p  �x�C�D98tA�� �M;�u���  �������@HQ�K�@,��ЋU����C�   �D��<����M��T�����l�����\������l�T�\�Y��Y��Y��X�<����Y�d����X�D����X��������X�L����Y��X���t����Y��Y�|����X�(��Y������Y�������   �������@HQ�K,�@,�Ћ�j �@Hh�  �s,��p  �   ��������Ћ�p  ���I�I�,��T��\�f(��Y�����f(��Y�����X�����f(��Y������Y�����X��X�����f(��Y�$����X������X�f(��Y�����Y�����X�f(��Y�,����Y�4����X��X�f֣�   �X�f֋   f֫  ���   �\cP��   �\SX��  �\K`��  f(��Y�   �Y�`  f(��Y�  �Y�  �X�(��Y�0  �X���   �Y��Y�(  �X���8  �Y��Y�@  �X��X��X�� tHtHu#W�f(�f(��W�f(�(��
W�f(�(����  ���  �Y����  f(��Y��  ��l����Y��Y��  �X����  �Y��Y��X����  �Y��X��X����  �Y��X����  �Y�f֛  f֓  �X�f֋   ���c  �E�9C$��  3��}�I �C�������R�@H�@,�Ћ�������P��l����   ������P��D  ��  ��  �@0�`��   �h �Y��Y��p(�}��Y��X��@H�Y��Y���X��@8�Y��E    �X��@P�Y��X��@@�Y��X��@X�C�Y| �X�t`3����$    ��Sf(ԋD�� �L0��D0��XT0�D0��X͍@�D�X�f��f�L�f�D��M�CA�M;Lu��E�@���E��}�;C$������  �{$ �E�    �~  3��u�	��$    ����`  �� �  H�z  H�5  �C��l�����R�@H�@,����   ��  ��0  �E���  �   ����������Y����f(��Y������M��Y�����X��  (��Y������X�(��Y�������X��  ��|����X���   �E��Y������L�����8  �X�(��Y�����X�(��Y������|����X�(��Y�$������M��X��E��Y�����M��Y�4�����t�����t���(��Y�����]��X�(��Y�$����X�(��Y�,�����t����X�(��Y�<�������`����X��E��Y�4�����`����E��U�(��Y�,����X�(��]��Y�L����Y�D����Y�T����Y�D����Y�<����Y�T����C�M�Xދ��XЋ@H�Xߋ@,��l���R�U��]��]��Y�L����X��X��]��Ћ�������P������   ������P��  ���  �@���  ���  f(��E��@0�Y��Y��p8�X �xP�hX���X��@H�Y��X��@ �E���@���f(��Y�(��Y��X`�X�(��Y��X��@(�E��Y���T����`@�X@�E��M�(��Y��X�(��Y��X��M����  �E��Y����  �E��@0�Y��  �]��X��@H�Y��X��E��Y��]��E��]�(��Y��  �X�(��Y��X��E��Y��]��E��M�(��Y��  �X�(��Y����  �X��E��M����  �Y��E��@0�Y��  �]��X��@H�Y��X��E��Y��]��E��]�(��Y��  �X�(��Y��X��E��Y��]��]��E��M�(��Y��  �X�(��Y��X����  �Y��M����  �]��X0�Y��  �U��X��XH�Y��X��]��Y��U����  �C�u�Y��| �Y��Y���   �Y�(  �X��Y��E�    �X��}��Y����   �Y�  �X��X���  �Y�@  �X��X���  �u��Y��Y��Y��]�3��S�mċD��`����Yl8�YD8��t����X�L����Yd8�� �X��E��YD8��X�|����X��E��YD8��X��E��YD8��D8�(��YU��X�(��YM��X�@����Ym��X�T����@�D�Xm�(��YE��X�(��YE��Ye��X��X��X�f���XM��X�f�L�f�l��M��CA�M�;L������  �C��l�����R�@H�@,����   ��  ��0  �E���  �   ����\�����Y�d���f(��Y�\����M��Y�|����X��  (��Y�\����X�(��Y�l������X��  �U��X���(  �E��Y�d�����T�����@  �X�(��Y�l����X�(��Y�t����]��X�(��Y��������M��X��E��Y�|����M��Y������E��U�(��Y�t����]��X�(��Y������X�(��Y������U��X�(��Y��������M��X��E��Y������]��E��U�(��Y������X�(��]��Y������Y������Y������Y������Y������Y������C�M�Xދ��XЋ@H�Xߋ@,��l���R�U��]��]��Y������X��X��]��Ћ���L���P��,����   ��L���P��1  ���  �@���  ���  f(��E��@0�Y��Y��p8�X �xP�hX���X��@H�Y��X��@ �E���@���f(��Y�(��Y��X`�X�(��Y��X��@(�E��Y���L����`@�X@��`�����`���(��Y��X�(��Y��X���`������  �E��Y����  �E��@0�Y��  �]��X��@H�Y��X��E��Y��]���|�����|���(��Y��  �X�(��Y��X��E��Y���|�����t�����t���(��Y��  �X�(��Y����  �X��E���t������  �Y��E��@0�Y��  �]��X��@H�Y��X��E��Y��]��E��]�(��Y��  �X�(��Y��X��E��Y��]��]��E��M�(��Y��  �X�(��Y��X����  �Y��M����  �]��X0�Y��  �U��X��XH�Y��X��]��Y��U����  �Y��Y��C�Xދu�Y�| ��   �Y�   �X��Y��E�    �]��]��Y���  �Y��   �X��X���8  �Y�  �X��X��]��V  �E��u��}��Y��Y��Y��E�3����S�m��D�E��Yl8�YD8�e��X�T����Yd8�� �X��E��YD8��Xe��X��E��YD8��X��E��YD8��D8�(��YU��X�(��Y�|����X�@����Y�t����X�L����@�D�X�`���(��YE��X��Xm��X��X�(��YE��Ye�f���X��X�f�L�f�l��M��CA�M�;L�����3  �C��l�����R�@H�@,����  ��   ��8  �E���  �   ����������Y�����f(��Y������M��Y������X��  (��Y������X�(��Y��������X��  �U��X���(  �E��Y�������t�����@  �X�(��Y������X�(��Y������]��X�(��Y��������M��X��E��Y������M��Y������E��U�(��Y������]��X�(��Y������X�(��Y������U��X�(��Y��������M��X��E��Y������]��E��U�(��Y������X�(��]��Y������Y������Y������Y������Y������Y������C�M�Xދ��XЋ@H�Xߋ@,��l���R�U��]��]��Y������X��X��]��Ћ�������P�������   ������P��  ���  ���  ���  f(��Y`f(��Y@0�X �p(�hX(��Y��X�f(��Y@H�Xx���X��@8�Y���T����` �Y����  �X`�X��@P�Y��X���@����`@(��Y����  �]��X�(��Y����  �X�(��Y@��L����E�(��Y@0�}��X��YX8(��Y@H�X�(��Y@ �}��X�(��Y��]��XP�Y��u��X��E��Y��u��p(�Y��X����  (��Yx�X����  �E����  �E��Y@0�X�(��Y@H�X��E��Y@8��`����E��}�(��Y@ �Y��X�(��Y��Y��X��E��Y��}��X����  (��Yx�X����  �E����  �E��Y@0�X�(��Y@H�X��E��Y@8�}���|�����|���(��Y@ �Y��X�(��Y��X��E��Y���|����X���  �Y�   �C�u�YՃ| �E�    �X��E����   �Y�   �X���  �Y�0  �X��  �E��}��u��Y��Y��Y��X�@����X�T���3��X�L����E�S�m��D�E��Yl8�YD8�e��X�t����Yd8�� �X��E��YD8��Xe��X��E��YD8��X��E��YD8��D8�(��Y�`����X�(��YM��Ym��X��XM�@�D�X�(��YE��X�(��Y�|����Ye�f���X��X�f�L�f�l��M��CA�M�;L�����E�@���E�u;C$�������l����CP�X�  ���}��E�f�E���  �XCXf�E���   �XC`f�E���C ǅ\���������B  �}�j h% �C  �u��������P��8���P��0���P��蝞  ��������轞  ���  3�9s$t03��	��$    ����K���   ��@j j��F�;s$u�j ��B  �~E�f�CP�~E�f�CX�~E���f�C`�C �,B  ��h  P�[  ����   ��x  P���   �Ѝ�l  P�Z[  j h% �B  ������   j j �u����������������5��  ��_^[��]� ���Н  ��l  P�[  ��������3��t  _��^[��]� �Mj ��/  �����=�����h  P��Z  ����   ��x  P���   �Ѝ�l  P�Z  ��������3��  _��^[��]� �����VW��3�9~$t S3ۋ��F���P�  G����;~$u�[�FP�F$    ��  ��d  P�9Z  ǆp      ����   �F P���   �Ѓ�_^���U���VWh`bhd  h<h�  �/  ����t���a������3���M�@Q�@�Сj �@j��@�M�h�bQ�Ѓ��E�P�M���  �0Whu'  �T�  ��PVj ht'  �C�  ��PhN� 赝  ���M����  ��E�IP�I�у���_^��]��������������bW�f�	f�Af�I0f�IHf�If�I f�A8f�IPf�If�I(f�I@f�AX����������U����   �M�qX�I8�y(�A@�YAP�Y�f(��YQP�E��M��\��A �E��Y�f(��U��Q �YQ@�\��E�(��YA8�U��M��}��E�(��Q0�\��A�Y��Y�W��]��e��X��AH�Y��X���bf.џ��DzB�Ef�f�@f�H0f�HHf�Hf�H f�@8f�HPf�Hf�H(f�H@f�@X��]��^��y�E��A(��Y�(��Yq@(��Ya8�(��YYP(��Yy �\��e�(��\��e��YA0�\e��YIH�\u��\��i�X��E��\E��Y��Y��Y��Y�V�X�W�YM���8����I�YM�(��\��\��YAH�Yy0�X��X��]��Y���@����E��\E��Y��QH(��YI@�X��E��Y��X��y0��P����E��Y��Y���X����E��Y���H�����`���(��YAX�\�(��YA(�Y���h���(��YIX�\��Y���p���(��YA@(��YI(�E��8������\�(��YA8�YU��Y���x���(��YIP�Y}��\�(��Yi8�YAP�Y��\��\й   �M��Y��Y��m��U��_^��]��U��V�@�u�@V�СV�@�u�@�С���@�΋@<�Ћj��Qj��u�RLP���ҋ�^]������������U��V����a���������  �Et	V�|  ����^]� ��U����`�@HV�@,W�U�R�Ћ��E�   ���_^��]� ̡j �@Hh�  ��p  Q�Ѓ������U��V�@�u�@V�Ћj �Ij��IhHbV�у���^]� ��������̸N� �����������U�����@h�u�@,Q�M�Q�ЋM�~ f��~@f�A�~@��f�A����]� �����������U����X���   ���E�Pǁ�    f �?  �����  ��MЋ@V�@Q�Сj �@j��@�M�hHcQ�С�u��@�M��@(Q�Ћ���I�E��IP�ы�A�M��@QV�С�M��@Q�@�С�M��@Q�@�С�M��@Q�@�M�Q�С��8�@�M��@<�Ћj��Qj��M�QP�BL�M��ЍE�P�7  ��M��@Q�@�С�M��@Q�@�С�MЋ@Q�@�Ѓ�^������]������������������������U��E��PV=�  ��  t+�� tH�T  ����  �����^��]ø   ^��]ËE3�90�(  SW�@�<�����^  �lc�Ȋ:u��t�Y:Zu������u�3��Ƀ�����   �tc�ȍd$ �:u��t�Y:Zu������u�3��Ƀ�����   ��c�Ȋ:u��t�Y:Zu������u�3��Ƀ���u;���M��@Q�@�Сj �@j��@�M�h�cQ�ЍE�P�]5  �M��v��c�I �:u��t�P:Qu������u�3�������uV��    �  �H��M��@Q�@�Сj �@j��@�M�h|cQ�ЍE�P��4  �M�Q�@�@�Ѓ��EF;0�����_[3�^��]�=�  ��   �u����   �~ ��   ��MЋ@Q�@�Сj �@j��@�M�h�cQ�Ћ���E�P�c�  P�E�P�E�P�����P�O4  ��M��@Q�@�С�M��@Q�@�С�MЋ@Q�@�Ѓ�3�^��]���U�����t]��]����������������U���E��t�I�   ;�j B�j P���   �Ѓ�]ù   ;�VB�W�xW�* ������u_^]�Wj V�+ �������_�F��   ^]�������������U��M��t+�=� t�y���A�u	�E]��) ��@�M� ]��]����������U��M��t+�=� t�y���A�u	�E]�) ��@�M� ]��]����������U���E��t�I�   ;�j B�j P���   �Ѓ�]ù   ;�VB�W�xW�) ������u_^]�Wj V�* �������_�F��   ^]�������������U���E��t�I�   ;�j B�j P���   �Ѓ�]ù   ;�VB�W�xW�) ������u_^]�Wj V�) �������_�F��   ^]�������������U���E��t�I�   ;�j B�j P���   �Ѓ�]ù   ;�VB�W�xW�( ������u_^]�Wj V�) �������_�F��   ^]�������������U���u�@� �Ѓ�]����������U���u�@� �Ѓ�]����������U��M��t��@�M��@  ]��]áhﾭދ@��@  ��Y����������U��V�u���t�Q�@� �Ѓ��    ^]�����������U���@���  ]��������������U��E��t�x��u�   ]�3�]������U���@��  ]�������������̡�@��   ��U���E��t!�u�I�u�   ;�B�P���   �Ѓ�]ù   ;�VB�W�xW��& ������u_^]�Wj V�d' �������_�F��   ^]�����������U��M��ɺ   Dʅ�t�u�@�u���   Q�Ѓ�]Ã�VB�W�yW�k& ������u_^]�Wj V��& �������_�F��   ^]����������������U���u�@� �Ѓ�]����������U���u�@� �Ѓ�]����������U��E�   ;�VB�W�xW��% ������u_^]Ã} tWj V�I& ��_������F��   ^]����������������U���E��t;�} �u�I�u�   t;�B�P���   �Ѓ�]Ã�B�P���  �Ѓ�]ù   ;�VB�W�xW�,% ������u_^]Ã} tWj V�% ��_������F��   ^]�����������U��M��ɺ   Dʅ�t*�} �u�@�uQt���   �Ѓ�]Ë��  �Ѓ�]Ã�VB�W�yW�$ ������u_^]�Wj V�% �������_�F��   ^]�������������U���u�@� �Ѓ�]����������U���u�@� �Ѓ�]������������c������������c���������̅�t�j������̡�@��  ���@��(  ��U�����@�U䋀   R�ЋMP���  �M��5�  �E��]� �����������̡�@��$  ��U���@��  ]��������������U���@���  ]�������������̡�@��  ��U���@���  ]��������������U���@��x  ]��������������U���@��|  ]�������������̡�@��d  ��U���@��p  ]��������������U���@��t  ]��������������U���EV����ct	V��������^]� �������������̡V�@j �@j����Ћ�^���������U��V�@j �u�@���Ћ�^]� �U��V�@�u�@j����Ћ�^]� ̡�@�@�����U��V�@j ���   ��Mj V�Ћ�^]� �����������U���u�@Q�@�Ѓ�]� �����U���u�@Q�@�Ѓ����@]� U��h#  �u�@�u�@l��]� �U��hF  �u�@�u�@l��]� �U���u�@�@t�ЋP���   �@X�Ѓ�]� ����U���u�@�@t�Ћ�u�Ћ��   R�@`�Ѓ�]� ���������������U���u�@���   �Ћȅ�u]� �Q���   �@�Ѓ�]� ��������U���@���   ]�������������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������3�� �����������3�� �����������U��M�E�A4�E�A �E��E�A0�E�A�l �A8 �A<# �A@�s �AD( �AH2 �AL- �AP�s �Al�s �AX�s �A\�s �A`A �Ad< �AT�s �Ah7 �Ap�s �At�s �A(�A,    ]��������������U���   h�   ��`���j P�$ j �u��`����u�u�uP�����E h�   �E���`���P�u�uj�K'  ��8��]�����U���   V�����  �����   S�u�M��9�  ��M��@Q�@�Сj �@j��@�M�hdQ�Ѓ��E�P�M����  j j��E�P�E�P��d���P�7�  ��P�E�P�:�  ��P�E�P�-�  ���P���  ���M����4�  �M��,�  ��d����!�  �M���  ��M��@Q�@�Ѓ��M����  ��[t	V��  ����^��]� ������U��V�u����  �����^]� ������Q���  YË�`��` ��`$��`,��`0��`<��`@��`�Q�@L���   �Ѓ�������������U���u�@L�u���   Q�Ѓ�]� ���������������U��V�@L�񋀠   V�Ћȡ����u�@LQ�u���   V�Ѓ�^]� ���   �@P�ЋP���   �M�BH��^]� �������������̡Q�@L��(  �Ѓ�������������U���u�@L�u��,  Q�Ѓ�]� ��������������̡�@L� ������U��V�@@�u�@�6�Ѓ��    ^]��������������̡�@L���   ��U��V�@@�u�@�6�Ѓ��    ^]���������������U�����@L�u�@Q�M�Q�ЋM��P�9����M��Q����E��]� ��������U���u�@L�u�@Q�Ѓ�]� ��U���u�@LQ���   �Ѓ�]� �̡Q�@L�@�Ѓ���������������̡Q�@L�@�Ѓ���������������̡Q�@L�@�Ѓ����������������U���u��u�@L�u�@ Q�Ѓ�]� ���������������U���u�@LQ��4  �Ѓ�]� ��U���u��u�@L�u�@$Q�Ѓ�]� ���������������U���u��u�@L�u�@(�uQ�Ѓ�]� �����������̡Q�@L�@,�Ѓ���������������̡Q�@L�@0�Ѓ���������������̡Q�@L�@4�Ѓ���������������̡j �@LQ�@8�Ѓ��������������U���u�@L�u��  Q�Ѓ�]� ���������������U���@L���   ]��������������U���@L���   ]��������������U���@L��l  ]��������������U���@L���   ]��������������U���@L���   ]��������������U���@L���   ]��������������U���@L���   ]��������������U���@L���   ]��������������U���@L���   ]��������������U���u�@LQ�@<�Ѓ�]� �����U���@L���   ]�������������̡Q�@L�@��Y�U���u�@L�u�@@Q�Ѓ�]� ��U��j �@L�u�@DQ�Ѓ�]� ���U��j�@L�u�@DQ�Ѓ�]� ���U��j �@L�u�@HQ�Ѓ�]� ���U��j�@L�u�@HQ�Ѓ�]� ��̡Q�@L���   �Ѓ�������������U�����@L�u��  Q�M�Q�ЋM��P������M�������E��]� �����U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    ��  j �E�P�E�P����  ���M����y�  ��t3����M܋��   Q�@8�Ѓ�����E܋��   P�	�у���^[��]����������U���$V�E��P�M��E�   �E�   �E��  �E�    �E�    �h�  j�E�P�E�P���7�  �M��ߌ  ��M܋��   Q� �Ѓ�^��]�����U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    ���  j �E�P�E�P����  ���M����i�  ��t
�M��  � ��M܋��   Q�@L�ЋM��P�{�  ��E܋��   P�	�ыE��^[��]� ���������U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    �G�  j �E�P�E�P�����  ���M���蹋  ��t
�M�=�  � ��M܋��   Q�@L�ЋM��P�˜  ��E܋��   P�	�ыE��^[��]� ���������U���$�V�u�E�    �E�    ���   ��@(�M�Q�Ѓ��E�P�M��E��  �E�    �E�    �~�  j�E�P�E�P���M�  �M����  ��M܋��   Q� �Ѓ�^��]� ��������U���$�V�u�E�    �E�    ���   ��@(�M�Q�Ѓ��E�P�M��E��  �E�    �E�    ��  j�E�P�E�P����  �M��e�  ��M܋��   Q� �Ѓ�^��]� ��������U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    �w�  j �E�P�E�P���&�  ���M�����  ^��[tW��E��E����M܋��   Q�@<�Ѓ���]��M܋��   Q� ���E�����]����������������U����EV�E��P�M�E�   �E��E��  �E�    �E�    �Ň  j�E�P�EP����  �M�<�  ��M䋀�   Q� �Ѓ�^��]� ���������������U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    �G�  j �E�P�E�P�����  ���M���蹈  ��t3����M܋��   Q�@8�Ѓ�����E܋��   P�	�у���^[��]����������U���$�EV�E�E��P�M��E�   �E��  �E�    �E�    詆  j�E�P�E�P���x�  �M�� �  ��M܋��   Q� �Ѓ�^��]� ���U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    �7�  j �E�P�E�P�����  ���M���詇  ��t8��u���   W��	���b�E�P�F�у���^[��]� ��M܋��   Q�@P���~ �u�f��~@���   �E܋	Pf�F�у���^[��]� ���U���$�V�u�E�    �E�    ���   ��@,�M�Q�Ѓ��E�P�M��E��  �E�    �E�    �>�  j�E�P�E�P����  �M�赆  ��M܋��   Q� �Ѓ�^��]� ��������U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    �Ǆ  j �E�P�E�P���v�  ���M����9�  ��t8��u���   W��	���b�E�P�F�у���^[��]� ��M܋��   Q�@P���~ �u�f��~@���   �E܋	Pf�F�у���^[��]� ���U���$�V�u�E�    �E�    ���   ��@,�M�Q�Ѓ��E�P�M��E��  �E�    �E�    �΃  j�E�P�E�P����  �M��E�  ��M܋��   Q� �Ѓ�^��]� ��������U�����@Lj�u���   Q�M�Q�ЋM�~ f��~@��f�A����]� U�����@Lj �u���   Q�M�Q�ЋM�~ f��~@��f�A����]� U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    �ׂ  j �E�P�E�P����  ���M����I�  ��t8��u���   W��	���b�E�P�F�у���^[��]� ��M܋��   Q�@P���~ �u�f��~@���   �E܋	Pf�F�у���^[��]� ���U���$�V�u�E�    �E�    ���   ��@,�M�Q�Ѓ��E�P�M��E��  �E�    �E�    �ށ  j�E�P�E�P����  �M��U�  ��M܋��   Q� �Ѓ�^��]� ��������U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    �g�  j �E�P�E�P����  ���M����ق  ��t8��u���   W��	���b�E�P�F�у���^[��]� ��M܋��   Q�@P���~ �u�f��~@���   �E܋	Pf�F�у���^[��]� ���U���$�V�u�E�    �E�    ���   ��@,�M�Q�Ѓ��E�P�M��E��  �E�    �E�    �n�  j�E�P�E�P���=�  �M���  ��M܋��   Q� �Ѓ�^��]� ��������U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    ��  j �E�P�E�P����  ���M����i�  ��t3����M܋��   Q�@8�Ѓ�����E܋��   P�	�у���^[��]����������U���$�EV�E�E��P�M��E�   �E��  �E�    �E�    �Y  j�E�P�E�P���(�  �M��Ѐ  ��M܋��   Q� �Ѓ�^��]� ���U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    ��~  j �E�P�E�P����  ���M����Y�  ��t8��u���   W��	���b�E�P�F�у���^[��]� ��M܋��   Q�@P���~ �u�f��~@���   �E܋	Pf�F�у���^[��]� ���U���$�V�u�E�    �E�    ���   ��@,�M�Q�Ѓ��E�P�M��E��  �E�    �E�    ��}  j�E�P�E�P����  �M��e  ��M܋��   Q� �Ѓ�^��]� ��������U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    �w}  j �E�P�E�P���&�  ���M�����~  ��t3����M܋��   Q�@8�Ѓ�����E܋��   P�	�у���^[��]����������U���$�EV�E�E��P�M��E�   �E��  �E�    �E�    ��|  j�E�P�E�P����  �M��P~  ��M܋��   Q� �Ѓ�^��]� ���U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    �g|  j �E�P�E�P����  ���M�����}  ��t3����M܋��   Q�@8�Ѓ�����E܋��   P�	�у���^[��]����������U���$�EV�E�E��P�M��E�   �E��  �E�    �E�    ��{  h�   �E�P�E�P����  �M��=}  ��M܋��   Q� �Ѓ�^��]� �������t��t��t3�ø   ���̡Q�@L�@L�Ѓ���������������̡Q�@L�@P�Ѓ����������������U���u��u�@L�u���  Q�Ѓ�]� ������������U���u�@LQ��  �Ѓ�]� ��U���u�@LQ���   �Ѓ�]� �̡Q�@L�@X�Ѓ����������������U���u��u�@L�u�@\Q�Ѓ�]� ���������������U����0�@LS�@V���Ћ؅�u^[��]� W�M��r����u�E�Eء�E�    �E�    �E�    �E�    �E�    �]Ћ@h]  �@0�M��Сj ���   j �@S���Ѕ���   �S�@L�@�Ћ�������   �d$ ����   �΋R(�ҋ��E�Ph�   �u��*  ����tq�M��tj�j ���   ���   �ЋЅ�tO�V���   �ʋ@<�С�M苀�   Q���   �Ѓ���t�V�@@�@�Ѓ������d����*�S�@@�@�С�M苀�   Q���   �Ѓ�3ۍM���  �M��x���_^��[��]� ������������̡Q�@L�@`�Ѓ���������������̡Q�@L�@d�Ѓ����������������U���u�@LQ�@h�Ѓ�]� ����̡Q�@L��D  �Ѓ������������̡Q�@L�@l�Ѓ����������������U���u�@LQ���   �Ѓ�]� �̡�@L�@�����U��V�@@�u�@�6�Ѓ��    ^]��������������̡Q�@L���   ��Y�������������̡Q�@L���   �Ѓ�������������U���u��u�@L�u���   �u�uQ�Ѓ�]� ������U���u��u�@L�u���   Q�Ѓ�]� ������������U���u��u�@L�u��   �uQ�Ѓ�]� ���������U���u��u�@L�u��   Q�Ѓ�]� ������������U���@L��H  ]�������������̡�@L��L  ��U���@L��P  ]��������������U���@L��T  ]��������������U���@L��p  ]��������������U���@L��t  ]��������������U���@L���  ]��������������U���@L���  ]��������������U���@L���  ]�������������̡�@L���  ��U��U$V�u�Eh� h� h�� hД R�u �q�u�Q�u����@L�$�u���   VQ�Ѓ�4^]�  �������̡�@���   ���@���   ��U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U��V�@�u���   �6�Ѓ��    ^]������������U��V�@L�@�Ћ���u^]áj �u�@�u��h  �uV�Ѓ���u�V�@@�@�Ѓ�3���^]������������U��j �H�u�E�� P�u��h  �u�Ѓ�]�������U���@���   ]��������������U���@L���   ]��������������U���u ��u�@�u���   �u�u�u�u�Ѓ�]����U��� ��E�    �E�    �E�    �E�    �E�    �E�    �E�    ���   V���   �Ћu�E���t8��t4�j�QLP���   ���ЋE��E�E�Ph=���u��
  ������   ��M����   Q���   �Ѓ��M��E�    ��  ��^��]���������������U��� ��E�    �E�    �E�    �E�    �E�    �E�    �E�    ���   V���   �Ћu�E���t8��t4�j�QLP���   ���ЋE��E�E�Ph<���u���	  ������   ��M����   Q���   �Ѓ��M��E�    �  ��^��]���������������U���@L���   ]��������������U���@L���   ]�������������̡�@L��  ���@L��@  ��U��M�]� �����U��M�u��P]�U��M�u��u�P]��������������U���u�M�u��u�u�P]���������    �A    �A    �A    �A    �A    �A    ���������������̡���   �AP���   ��Y��������U���u�@8Q�@D�Ѓ�]� ����̡�@8�@<�����U��V�@8�u�@@�6�Ѓ��    ^]���������������U���u��u�@8�u�@�u�u�uQ�Ѓ�]� ������U���u��u�@8�u�@�u�uQ�Ѓ�]� ��������̡�@8� ������U��V�@8�u�@�6�Ѓ��    ^]���������������U���u��u�@8�u�@Q�Ѓ�]� ���������������U���u�@8�u�@Q�Ѓ�]� �̡Q�@8�@�Ѓ����������������U���u�@8Q�@ �Ѓ�]� �����U���u��u�@8�u�@$�u�uQ�Ѓ�]� ���������U���u�@8�u�@(Q�Ѓ�]� ��U���u��u�@8�u�@,Q�Ѓ�]� ���������������U���u��u�@8�u�@Q�Ѓ�]� ���������������U���u�@8�u�@0Q�Ѓ�]� ��U���u��u�@8�u�@4Q�Ѓ�]� ���������������U���u�@8Q�@8�Ѓ�]� �����U��M��P�APP�A@P�A0P�A P�AP���   Q�u�Ѓ�]�������������̡�@���   ���@���  ��U���@�@,]�����������������U���@���  ]��������������U��V�H�u�IV�ыV�I�I8�у���^]����̡�@�@<�����U���@�@@]����������������̡�@�@D����̡�@�@H�����U���@�@L]�����������������U���@�@P]�����������������U���@��<  ]��������������U���@��,  ]��������������U���u��u�@�u���   �u�uh�6  �Ѓ�]�����U���@�@]�����������������U���� �@�M��@Q�Сj �@j��@�M�h�dQ�С�M��@Q�@�С�M��@Q�@�M�Q�С�� �@�M��@<�Ћj��Qj��u�M�P�BL�С�M��@Q�@�С�M��@Q�@�С�M��@Q�@�Ѓ���]����U���@���  ]��������������U���@��8  ]��������������U�����@V��  �M�WQ�Ћ�}�IW�I���ыW�IV�I�ы�E��IP�I�у���_^��]����U�����@V��  �M�WQ�Ћ�}�IW�I���ыW�IV�I�ы�E��IP�I�у���_^��]����U���@��x  ]��������������U���@��|  ]��������������U���@���  ]��������������U���@���  ]��������������U���@���  ]��������������U���@�@T]�����������������U���@�@X]�����������������U���@�@\]����������������̡�@�@`�����U���@���  ]�������������̡�@�@d����̡�@�@h�����U���@�@l]�����������������U���@�@p]�����������������U���@�@t]�����������������U���@��D  ]��������������U���@��  ]��������������U���@�@x]�����������������U���@��@  ]��������������U��V�u���bz  �V�I�u�I|�у���^]���������U���@���   ]��������������U���@��d  ]��������������U���@��h  ]��������������U���@���  ]�������������̡�@���   ��U��V�u�������V�I���   �у���^]��������̡�@��`  ��U���@��  ]��������������U�����@�u���   �M�Q�ЋM�~ f��~@f�A�~@��f�A����]������������U���@���  ]��������������U���u�E����@�D$�E���   �$�u�Ѓ�]�����������U���@���   ]��������������U���@���   ]��������������U���@���  ]��������������U���@���  ]��������������U���@��   ]��������������U���@��  ]��������������U���@��l  ]�������������̡�@���  ��U���@���  ]��������������U���@���  ]��������������U���@���  ]��������������U���@���  ]��������������U���@���  ]��������������U�����@V���  W�u�M�Q�Ћ�}�IW�I���ыW�IV�I�ы�E��IP�I�у���_^��]�U�����@V���  W�u�M�Q�Ћ�}�IW�I���ыW�IV�I�ы�E��IP�I�у���_^��]�U���@���  ]��������������U���@���  ]��������������U�����U��@R���   �U�R�U�RQ�Ѓ����#E���]����������������U�����U��@R���   �U�R�U�RQ�Ѓ����#E���]����������������U�����U��@R���   �U�R�U�RQ�Ѓ����#E���]����������������U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U���@��  ]��������������U���@��\  ]��������������U�����H�u��t  �u�E�P�у����u  �M��u  �E��]��������U���@��H  ]��������������U���@��T  ]�������������̡�@��p  ��U���@��8  ]��������������U���  �� 3ŉE��EP�u������h   P��) ����x	=�  |#��h8d�@hH  ��0  �Ѓ��E� ��������@Q��4  h�d�ЋM�3̓���  ��]������������������������U���u(�E�u$�P�u ��u�@0�u���   �u�u�uRQ�Ѓ�(]�$ ������U���u(�E�u$�P�u ��u�@0�u���   �u�u�uRQ�Ѓ�(]�$ ������U���u(��u$�@0�u ���   �u�u�u�u�u�uQ�Ѓ�(]�$ ���������̡Q�@0���   �Ѓ�������������U���u�@0�u���   Q�Ѓ�]� ���������������U���u��u�@0�u���   �uQ�Ѓ�]� ��������̡Q�@0���   �Ѓ�������������U���u��u�@0�u���   �uQ�Ѓ�]� ��������̡�@0���   ��U��V�@0�u���   �6�Ѓ��    ^]������������U�����@V�u��X  �u�M��uQ�Ћuj �    �F    �P���   V�I�ы�E����   P�	�у� ��^��]����������U���4VhLGOg�M�������j �IP�E�hicMCP��X  �Ћ���E�    �E�    ���   j �@R�M�Q�С�M����   Q� �Ѓ� �M�������M����   Q�@T�Ѓ���u
�M�6���� ��M����   Q�@T�ЋM��P�T�����E����   P�	�ыE��^��]������U���@���  ]��������������U���@���  ]��������������U���@���  ]��������������U�����@V��t  Wj �u�M��u�u�uQ�Ћ�}�IW�I���ыW�IV�I�ы�E��IP�I�у�(��_^��]������U�����@V�u���  �u�M��u�uQ�Ћuj �    �F    �P���   V�I�ы�E����   P�	�у�$��^��]�������U����4�@��p  �Ѕ���   h���M�������u�@h���@4�M��С�u�@h���@4�M��Сj �@�M̋�X  Q�M�hicMCQ�Ћ���E�    �E�    ���   j �@R�M�Q�С�M����   Q� �С�M����   Q� �Ѓ�$�M��=�����]����������U����4�@V��p  �Ѕ�u��u�HV�I�у���^��]�Wh!���M�������u�@h!���@4�M��Сj �@�M̋�X  Q�M�hicMCQ�Ћ���E�    �E�    ���   j �@R�M�Q�С�M����   Q� �С�M����   Q�@H�Ћ�}�IW�I���ыW�AV�@�Ћ�E����   P�	�у�4�M��#�����_^��]������������U����4�@V��p  �Ѕ�u��u�HV�I�у���^��]�Wh����M�������u�@h����@4�M��Сj �@�M̋�X  Q�M�hicMCQ�Ћ���E�    �E�    ���   j �@R�M�Q�С�M����   Q� �С�M����   Q�@H�Ћ�}�IW�I���ыW�AV�@�Ћ�E����   P�	�у�4�M�������_^��]������������U����4�@��p  �Ѕ�u��]�Vh#���M�������u�@h#���@4�M��Сj �@�M̋�X  Q�M�hicMCQ�Ћ���E�    �E�    ���   j �@R�M�Q�С�M����   Q� �С�M����   Q�@8�Ћ�����   �E��	P�у�(�M�������^��]�������U����4�@��p  �Ѕ�u��]�Vhs���M�������u�@hs���@4�M��Сj �@�M̋�X  Q�M�hicMCQ�Ћ���E�    �E�    ���   j �@R�M�Q�С�M����   Q� �С�M����   Q�@8�Ћ�����   �E��	P�у�(�M��=�����^��]�������U���@���  ]��������������U���@���  ]��������������U���@��@  ]��������������U��V�u���t�Q�@��D  �Ѓ��    ^]�������U���@��H  ]��������������U���@��L  ]��������������U���@��P  ]��������������U���@��T  ]��������������U���@��X  ]��������������U���@��\  ]�������������̡�@��d  ��U���@��h  ]��������������U���@��l  ]��������������U���@���  ]�������������̡�@���  ��U���@���  ]�������������̡�@��P  ���@���  ��U�����@�u���  �M�Q�ЋM��P�׽���M������E��]���������U���@���  ]��������������U���@���  ]��������������U���@���  ]��������������U���@���  ]��������������U���@���  ]��������������U���@���  ]��������������U���@��l  ]��������������U���@���  ]��������������U���@���  ]��������������U���@��$  ]��������������U���@��(  ]��������������U���@��,  ]�������������̡�@��0  ���@��<  ��U���@��  ]��������������U���@��`  ]��������������U���@��\  ]��������������U���@d�@P]�����������������U��M�9 t��@d�M�@T]��]���U���u��u�@h�u� �uQ�Ѓ�]� �������������U���u��u�@h�u���   �uQ�Ѓ�]� ���������U���u��u�@h�u�@Q�Ѓ�]� ���������������U���u��u�@h�u�@ �u�uQ�Ѓ�]� ���������U���u��E�@h�����   �$Q�Ѓ�]� �����U���u��E�@h�����   �$Q�Ѓ�]� �����U���u�@h�u���   Q�Ѓ�]� ���������������U���u�@h�u���   Q�Ѓ�]� ���������������U���E����@h�u(���   �u$���D$�E�$�u�uQ�M�Q�ЋM�~ f��~@f�A�~@��(f�A����]�$ �������U���E����@h�u$���   ���D$�E�$�u�uQ�M�Q�ЋM�~ f��~@f�A�~@��$f�A����]�  ����������U����EVW�}�E�E��P�M��    �G    �E�    �E�    �vP  j W�E�P���(�  �M���Q  ��_^��]� ������U���u��u�@h�u���   �uQ�Ѓ�]� ���������U���u�@hQ���   �Ѓ�]� �̡�@h�@X�����U��M�9 t��@h�M�@\]��]���U���@h���   ]��������������U���@h���   ]��������������U���@h���   ]��������������U���u ��u�@h�u�@`�u�u�u�uQ�Ѓ� ]� ���U���u ��u�@h�u�@d�u�u�u�uQ�Ѓ� ]� ���U���u�@h�u�@hQ�Ѓ�]� ��U���u�@h�u�@lQ�Ѓ�]� ��U���u�@h�u�@pQ�Ѓ�]� ��U���u ��u�@h�u���   �u�u�u�uQ�Ѓ� ]� U���u ��u�@h�u���   �u�u�u�uQ�Ѓ� ]� U���u ��u�@h�u���   �u�u�u�uQ�Ѓ� ]� U���u��u�@h�u���   �u�uQ�Ѓ�]� ������U���u��u�@h�u���   �uQ�Ѓ�]� ���������U���u��u�@h�u�@tQ�Ѓ�]� ���������������U���u�@hQ�@x�Ѓ�]� �����U���@h���   ]��������������U���u��u�@h�u�@|Q�Ѓ�]� ���������������U���u �E����@h�D$�E���   �D$�E�$Q�Ѓ� ]� ���������������U���E�@H���@�$Q�Ѓ�]� ����������̡j �@HQ���   �Ѓ�����������U���u�@Hj ���   Q�Ѓ�]� �j�@HQ���   �Ѓ�����������U���u�@Hj���   Q�Ѓ�]� �j�@HQ���   �Ѓ����������U���u�@Hj���   Q�Ѓ�]� �Q�@H���  �Ѓ�������������U���u�@HQ���  �Ѓ�]� ��U���u�@HQ���  �Ѓ�]� ��U���u�@HQ���  �Ѓ�]� ��U���u�@H�u��  Q�Ѓ�]� ���������������U���u�@H�u��  Q�Ѓ�]� ��������������̡Q�@H���   �Ѓ�������������U��VW�u���ў  ������t��u�AHV���   W�Ѓ���_^]� �������U��VW�u���u�^�  ������t��u�AHV���   W�Ѓ���_^]� ����U���u�@H�u���   Q�Ѓ�]� ���������������U���u�@H�u���   Q�Ѓ�]� ���������������U���u�@HQ���   �Ѓ�]� �̡Q�@H���  �Ѓ�������������U���u��u�@H�u���  �u�uQ�Ѓ�]� ������U�����@HW���   j ��h�  W�Ѓ��} u�   _��]� Vh�  �O�  ��������   �j �IHV���   W�у��M��R�����u�@h�  �@0�M��С�E�@���@,�$h�  �M��Сj �@@�M�@(QV�Ѓ��M��Y���^�   _��]� ^3�_��]� �̡Q�@H���   ��Y��������������U���u�@HQ���  �Ѓ�]� ��U���u�@HQ���  �Ѓ�]� �̡Q�@H��4  �Ѓ�������������U���@H� ]��U��V�@@�u�@�6�Ѓ��    ^]���������������U��S�]V�uW�> ��u3�S�@HW���   �Ѓ���u�j�@HW���   �Ѓ���t�   ��u����   �W�@H���   �Ѓ��} u!�u��u�@H�u���  VSW�Ѓ��I�ΉM��t@�u��u�V�u�@HQ���  SW�С�M���   ���@(�ЋȉE��uǋu�E�8 u�W�@H���   �Ѓ���t3���   �EW���@H��u$���   �СS�@HW���   �Ѓ�_^[]� ���   �С���} �@Hu�u���  j �uVSW�Ѓ�_^[]� � h  �Ѓ��E��u_^[]� ��΋��   �@x�ЋP���   �M�B|�Ѕ�tP�u�j �u�@HV���  SW�Ћȃ���t��u���   �@H�С�΋��   �@(�Ћ���u��E_^[]� U���u��u�@H�u���  �u�uQ�Ѓ�]� �����̡Q�@H���   ��Y�������������̡Q�@H���   �Ѓ�������������U���u�@H�u���   Q�Ѓ�]� ��������������̡Q�@H���   ��Y�������������̡Q�@H��t  ��Y�������������̡Q�@H��P  �Ѓ������������̡Q�@H��T  �Ѓ������������̡Q�@H��X  �Ѓ�������������U�����@HQ��\  �M�Q�ЋM�~ f��~@f�A�~@��f�A����]� ����������̡Q�@H��`  �Ѓ�������������U���u�@HQ��d  �Ѓ�]� ��U���E�@H����h  �$Q�Ѓ�]� ��������U���E�@H����t  �$Q�Ѓ�]� ��������U���E�@H����l  �$Q�Ѓ�]� ��������U���u�@HQ��p  �Ѓ�]� ��U���u��u�@H�u���  �uQ�Ѓ�]� ���������U���u��u�@H�u���  �u�u�uQ�Ѓ�]� ��̡h�  �@H� �Ѓ�������������U��V�@@�u�@�6�Ѓ��    ^]��������������̡Q�@H���   �Ѓ������������̡Q�@H���   �Ѓ�������������U���u�@HQ���   �Ѓ�]� ��U���u�@HQ���   �Ѓ�]� ��U���u�@H�u���  Q�Ѓ�]� ���������������U���u�@H�u��   Q�Ѓ�]� ���������������U���u��E�@H�����  �$Q�Ѓ�]� �����U��V�@Hh  � �Ћ�������   �uh�  �A�  �Ѓ���t^�j �AHR���   V���uh(  ��  �Ѓ���t3�j �AHR���   V�С�����   j �@j���Ћ�^]áV�@@�@�Ѓ�3�^]�����U��V�@@�u�@�6�Ѓ��    ^]��������������̡Q�@H��  �Ѓ������������̡Q�@H��  �Ѓ������������̡Q�@H���  �Ѓ������������̡Q�@H���  �Ѓ������������̡Q�@H���  �Ѓ�������������U���u�@H�u��  Q�Ѓ�]� ���������������U���u��u�@H�u��   Q�Ѓ�]� ������������U���u��u�@H�u��|  �uQ�Ѓ�]� ���������U��EV���u��@H���  �'��u��@H���  ���u(��@H���  V�Ѓ���tP�u���   ^]� 3�^]� ����������U���SW���   �؅���   �} ��   �V�AHj ��p  h�  W�Ћ���IHh�  ���   W�u��������E����   �u3��Ή}��  ����   �E�P�E�P�u��W��  ��t\�u�;u�T������u�U����ɋD�;D�t-��Hl����P�E�p�A�ЋD������tP���  F;u�~��}��MG�}��  �u;��v���^_��[��]� _3�[��]� U����V�@Hj ��p  ��h�  V�u��Ѓ��E���u^��]� �EW��u��@H���  �+��u��@H���  ����T  ��@H���  V�Ћ������6  S���O  �h�  �@H3ۋ��   V�]��Ѓ�����   �E����s�E��M�@lS�q�@�Ћ؃�����   ��s�I\�u�I,�у���t�F�P���v  ��s�@\�u�@,�Ѓ���t�F�P���Q  �M�;At"��s�@\�u�@,�Ѓ���tV���%  ��s�@\�u�@,�Ѓ���t�FP���   ��]��@H�E���   h�  �u�C�]����Ѓ�;�����[_�   ^��]� _3�^��]� ������̡Q�@H���  �Ѓ�������������U���u�@H�u���  Q�Ѓ�]� ���������������U���u��u�@H�u���  Q�Ѓ�]� �����������̡Q�@H���  �Ѓ������������̡Q�@H���  �Ѓ�������������U���u�@HQ��  �Ѓ�]� ��U���u�@HQ��  �Ѓ�]� �̡Q�@H��  �Ѓ�������������U���u�@HQ��  �Ѓ�]� �̡Q�@H��T  �Ѓ�������������U���u�@H�u��  Q�Ѓ�]� ���������������U���u�@HQ��8  �Ѓ�]� ��U���u�@HQ��<  �Ѓ�]� ��U���u��u�@H�u��@  Q�Ѓ�]� ������������U���u�@HQ���  �Ѓ�]� ��U���u�@HQ��H  �Ѓ�]� �̡Q�@H��L  ��Y��������������U��V�@Hh�  � �Ћ�����u^]á�u�@H�u��  V�Ѓ���u�V�@@�@�Ѓ�3���^]����������U��V�@@�u�@�6�Ѓ��    ^]���������������U���u��u�@H�u��   Q�Ѓ�]� ������������U���E�@H����$  �$Q�Ѓ�]� �������̡Q�@H��(  �Ѓ�������������U���u�@H�u��,  Q�Ѓ�]� ��������������̡�@H��  ��U���@H��  ]�������������̡V�@@��@,WV�Ћ���ȋBj ���   h�  �Ћh�  �IHV���   ���у���
��t_3�^Ë�_^�̡Q�@@�@,�Ћ���ЋAj ���   h�  �������U���E�@H����  �u�u���$Q�M�Q�ЋM�~ f��~@f�A�~@��f�A����]� ��������U���E�@H����  �u�u���$Q�M�Q�ЋM�~ f��~@f�A�~@��f�A����]� �������̡Q�@H���  �Ѓ�������������U���u�@H�u��8  Q�Ѓ�]� ���������������U���u��E�@H����0  �$�uQ�Ѓ�]� ��U���@H�@]�����������������U��V�@@�u�@�6�Ѓ��    ^]���������������U���u �E�u����@H�$�u���   �u�u�Ѓ�]�������������U���u�E����@H�$�u���   �u�u�Ѓ�]�����������������    ���������̡j�@H�1��|  �Ѓ����������U��V�@H�u��x  ����3Ƀ������^��]� ���̡j �@H�1��|  �Ѓ����������U��fnE�M����YE�Xe�,�;�}��]�;EOE]����������������U���H�S�@HV���   W�}h�  W�Ћ3��IHV���   ��h�  W�]��у��E��u�u��u����	  ��ϋ��   �@��=�  ���  �@HV���   h:  W�Ћh�  �IHW���   �E��ыV�IHh�  ���   W�E��u��ы�؋IHW��  �]��ыW�IH�E̋��  �у�(3��E�9u���   �C�E�3ۍ�$    �M̅�tNj�W�!�  ���t>�Mȍ@�|� ���M�~�� ��%�������;�u+蟤  �M�;�O��b�  ���E��M�� ;Au������E�G���E�;}�|��]ԋ]�E�}��tyj W����  ����  �M����  ��t[�M�蔇  �M�;�uL��I�@h�d���  ��h�  Q�M��Ѓ��EĉE���:  �M��p�  �u�P�u�褾  ���E�h�d�@����@h�  ���  Q�M��Ѓ��E�����  �u��u�P�`�  �Mԃ���~,�h�d�@�����   h�  Q�Ѓ��E����  �j��@HV��  W�Ѓ�����  �u��t jW�����  ���t  ���ˌ  ���E��3��uܡj �@Hh�  ���   W�ЉE�3�3҃��U��E�9E��  �{�}����    �M̅��/  j�P��  ����  �Mȍ@�|� �4��u�~�� ��%�������9E���  ���`�  3�3��E��E�    9^~|��������Шtf�E������������u�������L���E�T��N�E�L��E�J�L��N�E�L���E�J�L��N�E�uĉL���E�J�L��C;^|����  �Ǚ+�����~�M�QPQ�M��  �U��]��M܍R3��ÉE��+ÉEċƋ�;E���  �E���]���t5�E�U�[�]��~�f��~D�f�D�~D��ˋ]���f�D�E��U�[�~�f��~D�f�B�~D��ʋU�f�A;�}n�d$ �E�9�u_�L�����������w>�$��� �M�U�����-�M�U���T���M�U���T���M�U���T���U���;�|��M�E؃�B@�M�M܉U��E�;������;E���  �}��  �U���M�3�;G�Å���   �R�ƋG��@�~�f��~D�f�B�~D�f�B�G��@�E��~�f�B�~D�f�B �~D�f�B(��U��@�E��~ȍȍRf�D�0�~Af�D�8�~Af�D�@��t0�G�@�E��~ȍȍRf�D�H�~Af�D�P�~Af�D�X�G��u��@�E��~ȍȍRf���~Af�D��~Af�D��G��W��@�E�B�~ȍȍRf���~Af�D��~Af�D���W��@�E�B�~ȍȍRf���~Af�D��~Af�D��B�U���t8�G�@�E��~ȍȍRf���~Af�D��~Af�D��WB�U����G��}ЋU��Eԋu�@���Eԉ}�;E�������E�P菐���E�P膐������  �E�P�u����E�P�l����E�P�c�����3�_^[��]Ë��   �ϋ@��=  ��  �j �@Hh(  ���   W�Ћh(  �IHW���   ���у�3ɉEԅ�~���˅�t�|� �4Vu���A;�|�E�h�d�@����@hY  ���  Q�M��Ѓ��E�����   �u��u�P覸  �E�h�d��    �h^  �@Q���  �M��Ѓ��E��tD�u�SP�j�  ��ƋIH���   +���PVW�E��у���u�E�P�<����E�P�3�����_^3�[��]áj �@Hh�  ���   W�Ћj �IHh(  ���   W�E��ыȋE�3�3ۃ�3҉M��u��]؅��  �}䐋߅���   3��EЃ��~   �M��X�R�4v������I �E��E��~f��~Df�A�~Df�A�E�C�~Df�A�~D f�A �~D(�E�f�A(�}��;ǋEЍI0�v|��u��]؃|� tb�}�ƍ@�E��~ȍȍRBf���~Af�D��~Af�D��E��v�~ȍȍRBf���~Af�D��~Af�D��}�4ߋEԉu�C�]�;�������M��U�3���~#���$    ��    �D�    ��   @;�|�E�P胍�����E�P�w�����_^�   [��]�F� S� a� o� ��������U���u�E����@H�$�u���  �u�Ѓ�]���U���@H���  ]��������������U���@H���  ]��������������U���u0�E(����@H�$�u$���  �u �u�u�u�u�u�u�Ѓ�,]�U���@H���  ]��������������U���@H���  ]��������������U���u0�E�u,��u(�@H�u$��P  �u ���D$�E�$�u�u�Ѓ�,]��������������d�A    ����q��d��@l�@��Y���������U��V�@l��@�v�ЋM����u�A^]� �u��u�@lQ�u� ��3Ƀ������F^��]� �������������̋I��u3�áQ�@l�@�Ѓ������U�����U��@lR�@�U�R�u�u�q�ЋM��U��;�u	�E���]� ���9U�D���]� �������U���@H���   ]��������������U���@H���  ]��������������U�����M�@�����   W��$�u���]��E�M�f/�w�Ef/�w(���M�@���@,�$�u�Ћ�]����������U���0�W��M�Q�u�E��E��E��@�MЋ��   Q�M���~X�Ef/��~ �~P�Mv(��	f/�v(�f/�v(��	f/�v(�f/�wf/�v(��(ġ�E��U��]��@�M�@HQ�u�M�Ћ�]�������������U���@H��0  ]�������������̋������������������������������̡�@H���  ��U���@H���  ]��������������U���u0��u,�@H�u(���  �u$�u �u�u�u�u�u�uQ�Ѓ�0]�, ����U���u0��u,�@H�u(���  �u$�u �u�u�u�u�u�uQ�Ѓ�0]�, ���̡Q�@H��,  �Ѓ�������������U���u�@HQ��X  �Ѓ�]� �̡Q�@H��\  �Ѓ�������������U��Q�@H�u���   �u�Ѓ�]� ���������������U��QSV��MW�}3҉u��ϋ���t
����B��u��PSWV�M�	  �} ~(��   VW�}�W�M�o  SVW�M�  _^[��]� ;�tSWV�M�L  _^[��]� ���U��V���v��d��@l�@�Ѓ��Et	V���������^]� �����������U���V�u����   �ƙ+U��S��A�Z�W�	�<�ˉM��E��}�]���d$ �]��}�E���$    ��~I�����M��]��E��*�G���S����GN�C�u�}��W��~g�M��U����9u����    ���G���;�}��U;H}G���;�M��w������s��H�K�p�u�?��U;�~��M��N���_[^��]� �����U��UV�u��+����� ~^�E�U]�����S�ZW�]��I ��;�t7�]��$    �;H�}�p�ыH���H��H�P��p����;�u܋]�U�u���];�u�_[^]� ��U��QS�]W�}��+ǃ���M�=   ��   V�E��tu�7H�E��+����+����K��ǍǉU;�}9U|��;��;�}���9UL��M�PSW�u�   �u�M�S��V�u�z�����+������   �^_[��]� �M�SW�u�����^_[��]� ������������U��QS�]V�u;�t8W��F���;}$���N�M���
�H�@��J�R�;8|�E��:�B��;�u�_^[��]� U��ES�]VW�}�����9|���I ��;|�;�s$���p��O�H��w;�u����;�uǋ���_^[]� ���������̡Q�@\�@�Ѓ���������������̡Q�@\�@�Ѓ����������������U���u�@\Q�@�Ѓ�]� �����U���u�@\�u�@Q�Ѓ�]� ��U���u�@\Q�@�Ѓ�]� ����̡Q�@\�@�Ѓ����������������U���u�@\Q�@ �Ѓ�]� �����U���u�@\�u�@$Q�Ѓ�]� ��U���u��u�@\�u�@`�uQ�Ѓ�]� ������������U���u�@\Q�@0�Ѓ�]� �����U���u�@\Q�@@�Ѓ�]� �����U���u�@\Q�@D�Ѓ�]� �����U���u�@\Q�@H�Ѓ�]� ����̡Q�@\�@4�Ѓ����������������U���u�@\�u�@8Q�Ѓ�]� ��U���u�@\Q�@<�Ѓ�]� �����U���SVW�}��j �ω]��H  �S�@\�@�Ѓ���S���H  3���~?��I ��M��@\Q�@`�MQh���V�u��Ѓ����u�eH  �u����[H  F;�|�_^[��]� �������������U���S�]W�E��P���K  �}� |z�W�@\�@�Ѓ��E�P���K  �E���tWV3���~B�EP���}K  �E�P���rK  �M;M��Q�@\W�@�ЋMA���M;M�~�F;u�|�^_�   [��]� _�   [��]� ����������̡�@\� ������U��V�@\�u�@�6�Ѓ��    ^]����������������    �A    �A    �A    �����V��~ u=���t�Q�@<�@�Ѓ��    W�~��t����0  W�~�����F    _^���������U����E�VP���R  ����P�   �M���0  ��^��]���U��V��~ u4hej;h<j���������t�u���00  �3��F��u^]� �~ t3�9^��]� ��u�@<� �Ћȃ�3��ɉ�F   ��^]� �����V���F   ��@<�@��3Ʌ����^���������������U��	���u	�@� ]� �@<�u�@Q�Ѓ�]� �����̃y t�   ËQ��u3�áR�@<�1�@�Ѓ��������V��~ u=���t�Q�@<�@�Ѓ��    W�~��t���[/  W�u|�����F    _^���������U������u�@� ]Ë@<�u�@Q�Ѓ�]�������U�����$V��u��A�0���u�@<Q�@�Ћ�����I�E�ISP�ѡ�M�@Q�@V�С�M܋@Q�@�Сj �@j��@�M�h`eQ�С�� �@j �@@�M�Q�M�Q�M��Ѕ���M܋@Q�@���С����[t(�H�u�IV�ы�E�IP�I�у���^��]Ë@j�u��@H�M��Сj��@j��u�@L�u��M��С�u�@V�@�СV�H�E�IP�ы�E�IP�I�у���^��]������������U�����$SV��u��A�0���u�@<Q�@�Ћ�����I�E�IP�ѡ�M�@Q�@V�С�M܋@Q�@�Сj �@j��@�M�h`eQ�С�� �@j �@@�M�Q�M�Q�M��Ѕ���M܋@Q�@���С����t)�H�u�IV�ы�E�IP�I�у���^[��]Ë@j�u��@H�M��Сj��@j��u�@L�u��M��С�M܋@Q�@�Сj �@j��@�M�h`eQ�С���@j �@@�M�Q�M�Q�M��Ѕ���M܋@Q�@���С�����?����@j�u��@H�M��Сj��@j��u�@L�u��M��С�u�@V�@�СV�H�E�IP�ы�E�IP�I�у���^[��]���U�����$SV��u��A�0���u�@<Q�@�Ћ�����I�E�IP�ѡ�M�@Q�@V�С�M܋@Q�@�Сj �@j��@�M�h`eQ�С�� �@j �@@�M�Q�M�Q�M��Ѕ���M܋@Q�@���С����t)�H�u�IV�ы�E�IP�I�у���^[��]Ë@j�u��@H�M��Сj��@j��u�@L�u��M��С�M܋@Q�@�Сj �@j��@�M�h`eQ�С���@j �@@�M�Q�M�Q�M��Ѕ���M܋@Q�@���С�����?����@j�u��@H�M��Сj��@j��u�@L�u��M��С�M܋@Q�@�Сj �@j��@�M�h`eQ�С���@j �@@�M�Q�M�Q�M��Ѕ���M܋@Q�@���С����������@j�u��@H�M��Сj��@j��u�@L�u��M��С�u�@V�@�СV�H�E�IP�ы�E�IP�I�у���^[��]�����������U�����$SV��u��A�0���u�@<Q�@�Ћ�����I�E�IP�ѡ�M�@Q�@V�С�M܋@Q�@�Сj �@j��@�M�h`eQ�С�� �@j �@@�M�Q�M�Q�M��Ѕ���M܋@Q�@���С����t)�H�u�IV�ы�E�IP�I�у���^[��]Ë@j�u��@H�M��Сj��@j��u�@L�u��M��С�M܋@Q�@�Сj �@j��@�M�h`eQ�С���@j �@@�M�Q�M�Q�M��Ѕ���M܋@Q�@���С�����?����@j�u��@H�M��Сj��@j��u�@L�u��M��С�M܋@Q�@�Сj �@j��@�M�h`eQ�С���@j �@@�M�Q�M�Q�M��Ѕ���M܋@Q�@���С����������@j�u��@H�M��Сj��@j��u�@L�u��M��С�M܋@Q�@�Сj �@j��@�M�h`eQ�С���@j �@@�M�Q�M�Q�M��Ѕ���M܋@Q�@���С���������@j�u��@H�M��Сj��@j��u�@L�u��M��С�u�@V�@�СV�H�E�IP�ы�E�IP�I�у���^[��]���U��E����EȉM]�#  ������U���@<�@]�����������������U��E����u��]�VP�M��e�  �EP�E�P�M��E�    �E    藏  ����   �u�E���tA��t<��uX��u���   �@H�Ћ�ЋA���@xV���Ѕ�u+�   ^��]á�u���   �@T��VP�Y�������uՍEP�E�P�M���  ��u�3�^��]��������U���DS3ۉ]���M܋@V�@Q�СS�@j��@�M�hdeQ�С�M܋@<Q�@�Ћ���I�E܋IP�у���u^3�[��]�WV�M�3��9�  �E�P�E�P�M��y�  ���  ��}���   ��u����   �@T�Ћ�������   ����A�M̋@Q�С���@�M̋��   Qj�M�Q���Ћ���I�E܋IP�ы�A�M܋@QV�С�M��@Q�@�С���@�u�@x�M����E���t�E� ��t��M܋@Q�@����Ѓ���t��M̋@Q�@����Ѓ��}� u!�E�P�E�P�M��j�  ���������_^[��]Ë}���_^[��]��������������U���@SV�u3ۉ]���u^��M��@Q�@�СV�@j��@�M�hdeQ�С�M��@<Q�@�Ћ���I�E��IP�у���u^3�[��]�V�M��u�  �E�P�E�P�M�赌  ��t�W�}�E�����   ��u����   �@T�Ћ�������   ����A�MЋ@Q�С���@�MЋ��   Qj�M�Q���Ћ���I�E��IP�ы�A�M��@QV�С�M��@Q�@�С���@W�@x�M����E��t�E ��t��M��@Q�@����Ѓ���t��MЋ@Q�@����Ѓ��} tA�E�_^[��]Ã�u2�M���t+�Q���   �@H�Ћ�ЋA���@xW���Ѕ�t��E�P�E�P�M��f�  �������_^[��]�������̡�@<�@����̃=  uK����t�Q�@<�@�Ѓ���    V�5��t��� !  V�n�����    ^������������U���u��u�@�u���   �uQ�Ѓ�]� ���������U���u�E����@�D$�E���   �$�uQ�Ѓ�]� �������U���u��u�@�u���   Q�Ѓ�]� �����������̡Q�@���   �Ѓ�������������U���u��u�@�u���   Q�Ѓ�]� ������������U���u�@�u���   Q�Ѓ�]� ���������������U���u�@Q���  �Ѓ�]� ��U���u�@�@p�Ѓ�]� ������U���u�@�u���  Q�Ѓ�]� ���������������U���u�@�u���  Q�Ѓ�]� ���������������U���u�@�u���  Q�Ѓ�]� ���������������U���u�@�u���  Q�Ѓ�]� ���������������U����   V�u��u3�^��]�h�   ��0���j P蕖  ����M�Q���P��M��@�@<�Ѕ�tj �E�P�u�U�������u3���   �E��p����E��t����Eh�   ��0�����0���P�u��P����uǅ4����l j	�E��s �E��s �E�7 �E��s �E��s �E� �E�# ǅx����s ǅ|���( �E�< �E�A �E��s �E�F �E�K �E�P �E�U �E�Z �E�2 �E�- �E��s ����������E��IP�I�у���^��]�U��} u3�]� �W�u�P@����u_]� �w��u�@0�u���   �ЋG��_]� ���������U���u�@0�@�Ѓ���t��E   ��]�"]� ���̸   � ��������� ������������̃��� ����������� �������������U���u�H�I�ыE��]� ��̸   � ��������3�� ����������̸   @� ��������3��  ����������̸   � ��������3�� ��������������������������̸   � ��������3�� �����������3�� �����������U��E� ����]� �������������̸   � ��������U��E� ����]� ��������������3�� �����������U���@���  ]��������������U���@���  ]��������������U���   SV�u(W3�3��]����w  ��M�@�@<�Ѕ��F  �G  �E�����   �EP�M��n  ��M�@Q�@�СW�@j��@�M�hdQ�Ѓ��E�P�M��5  �u�Wj��E�P�E�P��\���P�_?�h<  ��P��x���P�h  ��P�E�P�[  ����P� C  �E���t�E� �� t�M�����S  ��t��x�������@  ��t��\�������-  ��t�M̃���  ��t��M�@Q�@����Ѓ���t�M���  �}� t�u(�u$�u��u�u�u���������E�P��E  ���V�u$j �u�u�u�����������E�IP�I�у���_^[��]��������������U���u�uj �u�u�u������]Ë�`��`��`��`��`��`(��`4��`8��`D��`H��`L��`P��`T�U��W�@j�@4���Mh�  ���u���u�F���_]� �U��V���PX�MP�  ��t�E^��   ]� �u���u�u�u�����^]� U��VW���Mj ��  �8�  �uuH� uB�j �@h�  ���   ���Ѕ�u�j �@h�  ���   ���Ѕ�t_3�^]� �u���u�u�uV�u�u���_^]� ���������������U���<S�]VW�}���`��u�F   WS�u���u�a���_^[��]� ����   j ���6  �8�  u8�i���P�F    �ܑ����M�@���@4jh�  ��_^�C�[��]� j ����  �8�  u�u��u���P_^�   [��]� j ����  �8�  tj ���  �8�G�����M�@j�@4h�  ���F    �$����������O�j	�PXP��j����3����U��E��t�P�IHR���  �у��E;F������~ �������M�@j ���   h�  �Ѕ�u"��M�@j ���   h�  �Ѕ��������M�@j �@4h�  �ЋM���t	j �x  ��E�F����   ���   �ЋM�E����   ����   Q聏�����M��֑���Mj�u�Yt���M�������E�E�E�E�E�ȉE��E�   �1�����t!HtHt	�E�    ��E�   ��E�   ��E�   �/����M���t�3����E�P����PXP�"����M�����t�3����M��{����M��s�����M���   Q���   �Ѓ��d�����M���   Q���   �Ѓ��   _^[��]� �������������A   �   � ��A   � ������U���u�A    ������]� �������U���u�@HQ���  �Ѓ�]� ��U��EV�0W�9;�t_3�^]� �P��u ��u9pu9qu��u�9yu�_�B^]� S�Y��u"��u9yu��u3��u/9pu*[_�   ^]� ��t��t;�u�P��t�A��t�;�t�[_3�^]� U���u�e������@]� ������������Vhj\hD ���~  ����t�@\��tV�Ѓ���^�����U��Vhj\hD ���Y~  ����t2�@\��t+V��hjxhD �7~  ����t�@x��t	V�u�Ѓ���^]� ���������U���Vhj\hD ����}  ����tG�@\��t@V�ЋEhjdhD �E��E�    �E�    ��}  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vhj\hD ���y}  ����t2�@\��t+V��hjdhD �W}  ����t�@d��t	�uV�Ѓ���^]� ���������U��Vhj\hD ���}  ����tZ�@\��tSV��hjdhD ��|  ����t�@d��t	�uV�Ѓ�hjhhD ��|  ����t�@h��t	�uV�Ѓ���^]� �U��Vhj\hD ���|  ������   �@\��t{V��hjdhD �s|  ����t�@d��t	�uV�Ѓ�hjhhD �K|  ����t�@h��t	�uV�Ѓ�hjhhD �#|  ����t�@h��t	�uV�Ѓ���^]� �����Vhj`hD ����{  ����t�@`��tV�Ѓ�^�������U��VhjdhD ���{  ����t�@d��t	�uV�Ѓ�^]� �������������U��VhjhhD ���y{  ����t�@h��t	�uV�Ѓ�^]� �������������VhjlhD ���<{  ����t�@l��tV�Ѓ�^�������U��VhjphD ���	{  ����t�@p��t�uV�Ѓ�^]� �^]� ���U��VhjxhD ����z  ����t�@x��t	V�u�Ѓ���^]� �����������U��Vhj|hD ���z  ����t�@|��tV�u�Ѓ�^]� 3�^]� ������U��Vhj|hD ���Iz  ����t�@|��tV�u�Ѓ����@^]� �   ^]� ��������������U���VhjthD ����y  ����tP�@t��tI�u�M�VQ�Ћu����P�`���hj`hD �y  ����th�H`��ta�E�P�у���^��]� hj\hD �y  �u����t4�@\��t-V��hjdhD �iy  ����t�@d��thV�Ѓ���^��]� �������U��Vhh�   hD ���&y  ����t���   ��t�uV�Ѓ�^]� 3�^]� U��Vhh�   hD ����x  ����t���   ��t�uV�Ѓ�^]� 3�^]� VW��3����$    �hjphD �x  ����t�@p��t	VW�Ѓ����8 tF��_��^�������U��SV��3�W��    hjphD �Ox  ����t�@p��t	VS�Ѓ����8 tphjphD �x  ����t�@p��tV�u�Ѓ�����hjphD ��w  ����t�@p��t	VS�Ѓ���W���x�����tF�^����E_��t�0��~=hjphD �w  ����t�@p��t	VS�Ѓ����8 u^�   []� ^3�[]� �����������U���Vhh�   hD ���Cw  ����t<���   ��t2�u�M�VQ��hj`hD �w  ����t�@`��t	�M�Q�Ѓ���^��]� �������U���Vhh�   hD ��v  ����tS���   ��tI�u�M��uQ�Ћu����P�:���hj`hD �v  ����td�H`��t]�E�P�у���^��]�hj\hD �jv  �u����t2�@\��t+V��hjxhD �Ev  ����t�@x��t	V�u�Ѓ���^��]�������̋���������������hjhD ��u  ����t	�@��t��3��������������U��V�u�> t+hjhD ��u  ����t�@��tV�Ѓ��    ^]�������U��} W��t0hjhD �u  ����t�@��t�u�uW�Ѓ�_]� 3�_]� �������������U��VhjhD ���9u  ����t�@��t�uV�Ѓ�^]� 3�^]� ������U��VhjhD ����t  ����t�@��t�uV�Ѓ�^]� 3�^]� ������Vhj hD ���t  ����t�@ ��tV�Ѓ�^�3�^���Vhj$hD ���t  ����t�@$��tV�Ѓ�^�3�^���U��Vhj(hD ���Yt  ����t�@(��t�u�u�uV�Ѓ�^]� 3�^]� U��Vhj,hD ���t  ����t�@,��t�u�uV�Ѓ�^]� 3�^]� ���U��Vhj(hD ����s  ����t�@0��t�u�u�uV�Ѓ�^]� 3�^]� Vhj4hD ���s  ����t�@4��tV�Ѓ�^�3�^���U��Vhj8hD ���is  ����t�@8��t�u�u�u�uV�Ѓ�^]� 3�^]� �������������U��Vhj<hD ���s  ����t�@<��t	�uV�Ѓ�^]� �������������U��Vhh�   hD ����r  ����u^]� �u���   V�Ѓ�^]� ������U��Vhh�   hD ���r  ����u^]� �u���   V�Ѓ�^]� ������U��Vhh�   hD ���Vr  ����u^]� �u���   V�Ѓ�^]� ������U��Vhh�   hD ���r  ����t�u���   �u�uV�Ѓ�^]� �����VhjDhD ����q  ����t�@D��tV�Ѓ�^�3�^���U��VhjHhD ���q  ����t�u�@HV�Ѓ�^]� �U��VhjLhD ���yq  ����u^]� �u�@LV�Ѓ�^]� ������������U��VhjPhD ���9q  ����u^]� �u�@P�uV�Ѓ�^]� ���������U��Vhh�   hD ����p  ����u^]� �u���   �u�uV�Ѓ�^]� U��Vhh�   hD ���p  ����u^]� �u���   �u�u�u�uV�Ѓ�^]� ����������VhjThD ���lp  ����u^Ë@TV�Ѓ�^���������U��VhjXhD ���9p  ����t�u�@XV�Ѓ�^]� �U���Vhh�   hD ���p  ����tQ���   ��tG�u�M�Q���ЋuP���l���hj`hD ��o  ����t|�H`��tu�E�P�у���^��]� hj\hD �E�    �E�    �E�    �o  �u����t3�@\��t,V��hjdhD �`o  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vhh�   hD ���o  ����t���   ��t�u���u�u��^]� 3�^]� ������������U��Vhh�   hD ����n  ����t���   ��t�u����^]� 3�^]� ��U��Vhh�   hD ���n  ����t���   ��t�u����^]� 3�^]� ��U��Vhh�   hD ���Fn  ����t���   ��t�u����^]� 3�^]� ��Vhh�   hD ���	n  ����t���   ��t��^��3�^����������������U��Vhh�   hD ����m  ����t���   ��t�u���u�u��^]� 3�^]� ������������U��Vhh�   hD ���vm  ����t���   ��t�u����^]� ���������U��Vhh�   hD ���6m  ����t���   ��t�u���u�u��^]� 3�^]� ������������Vhh�   hD ����l  ����t���   ��t��^��3�^����������������U��hjhD �l  ����t
�@��t]��3�]��������U���Vhh�   hD �ul  ����u��u�HV�I�у���^��]Ë��   W�u�M�Q�Ћ�}�IW�I���ыW�IV�I�ы�E��IP�I�у���_^��]���U��h�uhD ��k  ��]�������U��E�� ]�̡�@$�@X�����U���@$�@\]�����������������U���u��u�@$�u�@`Q�Ѓ�]� ��������������̡V�@��@V�СV�@$�@D�Ѓ���^�����������U��V�@��@V�СV�@$�@D�С�u�@$V�@d�Ѓ���^]� ���U��V�@��@V�СV�@$�@D�С�u�@$V�@�Ѓ���^]� ���U��V�@��@V�СV�@$�@D�СV�@$�u�@L�Ѓ���^]� ��̡V�@$��@HV�СV�@�@�Ѓ�^�������������U���u�@$Q�@L�Ѓ�]� �����U���@$�@]����������������̡Q�@$�@�Ѓ����������������U�����@$V�@WQ�M�Q�Ћ�}�IW�I���ыW�IV�I�ы�E��IP�I�у���_^��]� ���U���u�@$Q�@�Ѓ�]� �����U�����@$V�@ WQ�M�Q�Ћ�}�IW�I���ыW�A$�@D�СW�@$V�@L�С�H$�E�IHP�ы�E�IP�I�у� ��_^��]� ����U�����@$V�@$WQ�M�Q�Ћ�}�IW�I���ыW�A$�@D�СW�@$V�@L�С�H$�E�IHP�ы�E�IP�I�у� ��_^��]� ����U���,�E�VWP�o����P�I$�E�P�A�Ћ�}�IW�I���ыW�AV�@�С�M��@Q�@�С�H$�EԋIHP�ы�EԋIP�I�у� ��_^��]� ������̡Q�@$�@(��YáQ�@$�@h��Y�U���u�@$Q�@,�Ѓ�]� �����U���u�@$Q�@0�Ѓ�]� �����U���u�@$Q�@4�Ѓ�]� �����U���u�@$Q�@8�Ѓ�]� �����U���u�@$�u�@PQ�Ѓ�]� ��U���u�@$Q�@T�Ѓ�]� �����U���@$�@l]����������������̡�@$�@p�����U��V�@$��@LV�u�Ѓ���^]� ���������������U��V�@�u�@V�СV�@$�@D�СV�@$�u�@L�Ћ�u�I$V�I@�у���^]���U��V�@$�u�@@��V�Ѓ���^]� ���������������U���u�@$Q�@<�Ѓ�]� �����U���u�@$Q�@<�Ѓ����@]� U�����@$V�@tWQ�M�Q�Ћ�}�IW�I���ыW�IV�I�ы�E��IP�I�у���_^��]� ���U���@(�@]����������������̡�@(�@�����U���@(�@]�����������������U���@(�@]�����������������U���@(�@ ]�����������������U��j�u�@(�u�@��]� ����U���u��u�@(�u�@$��]� ��̡�@(�@(����̡�@(�@,����̡�@(�@0�����U���@(�@4]�����������������U���@(�@X]�����������������U���@(�@\]�����������������U���@(�@`]�����������������U���@(�@d]�����������������U���@(�@h]�����������������U���@(�@l]�����������������U���@(�@p]�����������������U���@(�@t]�����������������U���@(�@x]�����������������U���@(���   ]��������������U�����@V�@��M�Q�Ѓ��E�P���   ��u3����M��@$Q�u�@�Ѓ��   ��E��IP�I�у���^��]� ������U��Q��U��@(R�@X�Ѕ�u��]� �E3�8M�����   ��]� ���������U����V���E�    �E�    �@(�M��@hQ���Ѕ�t�M����u@�@�M�@Q�С�u�@�M�@Q�С�M�@Q�@�Ѓ��   ^��]� �@h�e���   hj  Q�Ћȡ���M��@(��u�@4j�����3�^��]� �@j �u�Q���Ѕ�u�E�P��F����3�^��]� �j �H�E�HP�u��A�u�ЍE�P�F�����   ^��]� ��U��V�@(W�}�@pW���Ѕ�t9��΋P(�GP�Bp�Ѕ�t"��΋P(�GP�Bp�Ѕ�t_�   ^]� _3�^]� ���U��V�@(W�}�@tW���Ѕ�t9��΋P(�GP�Bt�Ѕ�t"��΋P(�GP�Bt�Ѕ�t_�   ^]� _3�^]� ���U��S�@(V�@pW�}W���Ѕ���   ��΋P(�GP�Bp�Ѕ���   ��΋P(�GP�Bp�Ѕ�to��_�@(S�@p���Ѕ�tX��΋P(�CP�Bp�Ѕ�tA��΋P(�CP�Bp�Ѕ�t*�GP��������t�G$P��������t_^�   []� _^3�[]� �����U��S�@(V�@tW�}W���Ѕ���   ��΋P(�GP�Bt�Ѕ���   ��΋P(�GP�Bt�Ѕ�to��_�@(S�@t���Ѕ�tX��΋P(�CP�Bt�Ѕ�tA��΋P(�CP�Bt�Ѕ�t*�G0P���-�����t�GHP��������t_^�   []� _^3�[]� �����U���@(�@8]�����������������U���@(�@<]�����������������U���@(�@@]�����������������U���@(�@D]�����������������U���@(�@H]�����������������U���@(�@L]�����������������U���E�@(Q�@P�$��]� �U���E�@(���@T�$��]� ���������������U���u�@(�u�@|��]� ������U���u�@(�u���   ��]� ���U���� �@$V�@W�u���M�Q�Ћ���I�E��IP�ы�A�M��@QV�С�M��@Q�@�Ѓ��E�P���L   ����I�E��IP�у���_^��]� �����������U���} �P(�����E�B8]����U��Q�V�@W�@d���Mj �Ћh�e�I�p���   h�  V�ыȡ���M���u�@(j��@4����_3�^��]� �@j �@hVQ�M�СV�@(�ϋ@H�Ѕ�t�V�@(�u��@ ���Ѕ�t�   �3��E�P�tA������_^��]� �������U��V�@(W�}�@P�Q���$�Ѕ�tG��G�@(Q�@P���$�Ѕ�t)��G�@(Q�@P���$�Ѕ�t_�   ^]� _3�^]� ������������U��V�@(W�}�@T������$�Ѕ�tK��G�@(���@T���$�Ѕ�t+��G�@(���@T���$�Ѕ�t_�   ^]� _3�^]� ������U��V�@(W�}�@P�Q���$�Ѕ��  ��G�@(Q�@P���$�Ѕ���   ��G�@(Q�@P���$�Ѕ���   ��G�@(Q�@P���$�Ѕ���   ��G�@(Q�@P���$�Ѕ���   ��G�@(Q�@P���$�Ѕ�tt��G�@(Q�@P���$�Ѕ�tV��G�@(Q�@P���$�Ѕ�t8��G �@(Q�@P���$�Ѕ�t�G$P���������t_�   ^]� _3�^]� �����U��V�@(W�}�@T������$�Ѕ���   ��G�@(���@T���$�Ѕ���   ��G�@(���@T���$�Ѕ���   ��G�@(���@T���$�Ѕ�ti��G �@(���@T���$�Ѕ�tI��G(�@(���@T���$�Ѕ�t)�G0P���R�����t�GHP���C�����t_�   ^]� _3�^]� �����������̡�@(� ������U��V�@(�u�@�6�Ѓ��    ^]���������������U���@(���   ]��������������U���@(�@]����������������̡�@(�@�����U��V�@(�u�@�6�Ѓ��    ^]���������������U���u�@,�u�@Q�Ѓ�]� �̡�@,�@����̡�@,�@����̡�@,�@����̡�@,�@ ����̡�@,�@(����̡�@,�@$�����U���@,�@]�����������������U�����@,V�@W�U�R�Ћ�}�IW�I���ыW�A$�@D�СW�@$V�@L�С�H$�E�IHP�ы�E�IP�I�у���_^��]� ����̡j �@,j � �Ѓ��������������U��V�@,�u�@�6�Ѓ��    ^]��������������̡�@,�@4����̡�@,�@8�����U�����@,V�@<W�U�R�Ћ�}�IW�I���ыW�A$�@D�СW�@$V�@L�С�H$�E�IHP�ы�E�IP�I�у���_^��]� �����U�����@,V�@@W�u�U�R�Ћ�}�IW�I���ыW�IV�I�ы�E��IP�I�у���_^��]� ̡�@,�@,�����U��V�@,�u�@0�6�Ѓ��    ^]���������������U���@���  ]��������������U���@���  ]��������������U���@���  ]��������������U���@���  ]��������������U���@�@]�����������������U���@�@]�����������������U���@�@]�����������������U���@�@]�����������������U���@�@]�����������������U���@�@]�����������������U���u�@�u�@\��]� ������U���u�@�u��  ��]� ���U���E�@���@ �$��]� ���������������U���E�@Q�@$�$��]� �U���E�@���@(�$��]� ���������������U���@�@,]�����������������U���@�@0]�����������������U���@�@4]�����������������U���@�@8]�����������������U���@�@<]�����������������U���@�@@]�����������������U���@�@D]�����������������U���@�@H]�����������������U���@�@L]�����������������U���@�@P]�����������������U���@���   ]��������������U���u�@Q��  �Ѓ�]� ��U���@�@T]�����������������U���@�@X]�����������������U��U��u3�]� �R�@ Q�@(�Ѓ��   ]� �����U���@���   ]��������������U���@�@`]�����������������U���@�@d]�����������������U���@�@h]�����������������U���@�@l]�����������������U���@�@p]�����������������U���@�@t]�����������������U���@���   ]��������������U���@��  ]��������������U���@�@x]�����������������U���@�@|]�����������������U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U���u�@Q��  �Ѓ�]� ��U���@���   ]��������������U���@���   ]��������������U��U��t�R�@ Q�@$�Ѓ���t	�   ]� 3�]� �U��Q�@ �u�@L�u�Ѓ�]� ��U���@���   ]�������������̡�@���   ��U���@���   ]��������������U���@���   ]��������������U���@���   ]��������������U���@���   ]�������������̡�@���   ��U���@���   ]�������������̡�@���   ���@���   ���@���   ���@���   ���@���   ��U��V�@�u���   V�Ѓ��    ^]�������������U���@� ]���@�@�����U���@���   ]��������������U���@��   ]��������������U���@�@]�����������������U���@�@]�����������������U���@�@]�����������������U���@�@]�����������������U���@�@]�����������������U���@���  ]��������������U���@�@]�����������������U����E�V�uP���������M�@$Q�@�Ѓ���t]��M�@j�@Q�Ѓ���u�E�P��������t3�j�@V�@�Ѓ���u�V�@�@�Ѓ���t�   �3���H$�E�IHP�ы�E�IP�I�у���^��]��������U���@�@ ]�����������������U���@�@(]�����������������U���@��  ]��������������U���@��   ]��������������U���@��  ]��������������U���@��  ]��������������U�����@V�@$�M�WQ�Ћ�}�IW�I���ыW�A$�@D�СW�@$V�@L�С�H$�E�IHP�ы�E�IP�I�у���_^��]��������U�����@V���  �M�WQ�Ћ�}�IW�I���ыW�A$�@D�СW�@$V�@L�С�H$�E�IHP�ы�E�IP�I�у���_^��]�����U��j�u�  �E��]������������U���<�0SVW�E�    ��t�E�P�   �������-��M��@Q�@�   �С�M��@$Q�@D�Ѓ��}��u�@V�@�СV�@$�@D�СV�@$W�@L�Ѓ���t(��M��@$Q�@H����С�M��@Q�@�Ѓ���t&��H$�EċIHP�ы�EċIP�I�у�_��^[��]������U�����@V���  W�u�M�Q�Ћ�}�IW�I���ыW�A$�@D�СW�@$V�@L�С�H$�E�IHP�ы�E�IP�I�у� ��_^��]��U���@��D  ]��������������U���@��H  ]��������������U���@��L  ]��������������U�����@V���  W�u�M��uQ�Ћ�}�IW�I���ыW�IV�I�ы�E��IP�I�у���_^��]��������������U���@���  ]��������������U���@���  ]�������������̡�@��   ��U��V�@�u��$  �6�Ѓ��    ^]������������U��V�@��(  V�u�Ѓ���^]� ������������U��Q�@�u��,  �Ѓ�]� ��U��Q�@�u��,  �Ѓ����@]� �������������U��E��t�P�3ҡR�@Q��8  �Ѓ�]� ������U���u�@Q��<  �Ѓ�]� ��U���u��u�@�u��@  Q�Ѓ�]� ������������U���u�@�u��D  Q�Ѓ�]� ���������������U���u�@Q��H  �Ѓ�]� ��U�����@V��L  W�uQ�M�Q�Ћ�}�IW�I���ыW�IV�I�ы�E��IP�I�у���_^��]� ������������̡Q�@��T  �Ѓ������������̡Q�@��P  �Ѓ�������������U���u�@Q��X  �Ѓ�]� ��U���u�@Q��l  �Ѓ�]� �̡�@��0  ���@��4  ���@��p  ���@��t  ���@��\  ��U��V�@�u��`  �6�Ѓ��    ^]������������U���u��u�@�u��d  �u�uQ�Ѓ�]� ������U���u��u�@�u��h  �u�uQ�Ѓ�]� �����̡Q�@�@�Ѓ����������������U���u��u�@�u�@X�uQ�Ѓ�]� ������������U���u�@Q�@\�Ѓ�]� ����̡Q�@�@ ��Y�U�����@V���   h�  Q�M�Q�ЋP���   �@8�Ћ�����   �E��	P�у���^��]��������������U���@��   ]��������������U���u��u�@�u�@Q�Ѓ�]� ���������������U���u��u�@�u���   �uQ�Ѓ�]� ���������U���@�@$]�����������������U���u��u�@�u�@(�uQ�Ѓ�]� ������������U���u��u�@�u�@,�uQ�Ѓ�]� ������������U���u(��u$�@�u �@`�u�u�u�u�u�uQ�Ѓ�(]�$ �������������U��V�@W�@��W�ЋW�J���I���u��u�Q�u�N�QHP�B4j j W�Ѓ�(_^]� ���������������U���u ��u�@�u�@4�u�u�u�uQ�Ѓ� ]� ���U���u�@�u�@@Q�Ѓ�]� ��U���u�@Q�@D�Ѓ�]� ����̡Q�@�@L�Ѓ���������������̡Q�@�@L�Ѓ���������������̡Q�@�@P�Ѓ����������������U���u�@Q�@T�Ѓ�]� �����U���u�@Q�@T�Ѓ�]� ����̡Q�@�@h�Ѓ����������������U���u�@�u���   Q�Ѓ�]� ���������������U�����@V�u���   �uQ�M�Q�Ћuj �    �F    �P���   V�I�ы�E����   P�	�у� ��^��]� ��������̡�@� ������U��V�@�u�@�6�Ѓ��    ^]���������������U���u��u�@�u���   �u�uQ�Ѓ�]� ������U��V�@�u�@�6�Ѓ��    ^]���������������U��QS�]V�C    ���@V�@h�Ѓ����u"�@hXf��0  h�  �Ѓ�^3�[��]� �M�Q�MQ�u�E    �@V���   �Ѓ���t�3�9u�~*W��I �E�<� �<�tj����
  ��t��F;u�|�_�EP�S"�����   ^[��]� ���U��QS�]V�C    ���@V�@h�Ѓ����u"�@hXf��0  h�  �Ѓ�^3�[��]� �M�Q�MQ�u�E    �@V���   �Ѓ���tу} t�3�9u�~<W�E����t*�Q�@�@h�Ѓ���t�Ej�<����!
  ��t�8F;u�|�_�EP�{!�����   ^[��]� �����������U���@��x  ]�������������̡�@��|  ��Q�@���   �Ѓ�������������U���u�@Q���   �Ѓ�]� �̡�@���   ��U��V�@�u���   �6�Ѓ��    ^]������������VW���O����W�f�G f�G(f�G0f�G8f�G@f�GHf�GPf�GX�    �G`    �Gd    �Gh    �Gp�Gx�����G|   ��_^�������V���X   �N^�������������������W��    �A`    �Ad    �Ah    �Ap�Ax�����A|   ���������������SW�����t7���#���xP t$V���#��j j �pPj�GP���#���H ���^�    �O`��t�Q�@�@�Ѓ��G`    _[��������������hXfh�   h<h�   ��������t������3��������U��V�uW�>��t���K����O����W�����_�    ^]�U��S�@V��   W��W�_dS�wx�w`�uV�Ѓ��G|����   �? ��   �; ��   �wpV�_hS�u�P������u&�W���hXf�@h  ��0  �Ѓ��u�O��������W"���xP u����"���E"��j j �pPj�GP���1"���H ��ЉG|��t���[����G|_^[]� �G|�Gx����_^[]� �G|�����    ��6�@�@�Ѓ��    �G|_^[]� �V������W��    �F`    �Fd    �Fh    �Fp�Fx�����F|   ^������U��QW���d �G`t~S�];_xttV�7�ΉE�u��g!���xP u����#���U!���M�S�u�pPj�GP�@!���H ��ЉG|^��u�E�_x��t�    �G`[_��]� �M�Gx������t�3�[_��]� �����������U��E��t	�Ap� �yd t�Ah]� 3��y|��]� ���U���u ��u�@�u�@�u�u�u�uQ�Ѓ� ]� ���U���u�@Q�@�Ѓ�]� ����̡Q�@�@��Y�U���u�@�u�@Q�Ѓ�]� �̡�@� ������U��V�@�u�@�6�Ѓ��    ^]���������������U��VW�������u���u�x@�u�����H ���_^]� ����U��VW�������u���u�xD�u����H ���_^]� ����W������xH u3�_�V������ύpH�|���H �^_�����U��W���e���xL u3�_]� V���P���u���u�pL�u�=���H ���^_]� U��W���%���xP u���_]� V������u���u�pP�u�u�����H ���^_]� ������������U��W�������xT u���_]� V������u���u�pT����H ���^_]� ��U��W������xX u���_]� V������u�ύpX�r���H ���^_]� �����U���SVW�}�م�t.�M��������?���pL�E�P���1���H ��ЍM��  ���u��tW��M��@Q�@�С�M��@V�@Q�С�M��@Q�@�Ѓ��������H@��t�V�@Q�@�Ѓ�_^[��]� ���������U��VW������u�΍xH����H ���_^]� ����������U��W���u���x` u
� }  _]� V���]���u�ύp`�P���H ���^_]� ���U��SVW���3���x` u� }  �#������p`�E���P������H ��Ћ���]�IS�I�у�;�>�S�@�@�Ѓ�;�)�������u���u�pDS�u����H ���_^[]� _^�����[]� U��W������xP u
�����_]� V���}���u���u�pP�u�u�u�u�a���H ���^_]� ����U��W���E���xT u
�����_]� V���-���u���u�pT����H ���^_]� U��W������xX tV�������u�ύpX�����H ���^_]� �������������U����E�P�u�E�    �E�    �E�    �E�    �E�    �E�    ��4  ����t(�M��t!�u���u�@�u��@X�u�Q�Ѓ���]�3���]����������������U��USV��F�����N;�~}�W�@�+����ρ�  �yI���Au��u	�   +���h�f�Hh�   ��    P�6��  �ЋЃ���t�N�~_�^�^��[]� �F_�F^��[]� �^^[]� ���������������A    �    �A    �A   �����U���u��u�@@�u�@Q�Ѓ�]� ���������������U���u�@@Q�@�Ѓ�]� �����U���u�@@�u�@Q�Ѓ�]� ��U���u�@@Q�@ �Ѓ�]� �����U�����   �@]��������������U�����   �@]��������������U�����   �@ ]�������������̡���   �@$��U�����   ���   ]�����������U�����   ��D  ]�����������U���u�@@Q�@L�Ѓ�]� ����̡Q�@@�@H�Ѓ����������������U�����   ���   ]�����������U�����   ���   ]����������̡Q�@H���   �Ѓ�������������U��V��M��t2�U����   ��t�@@R��^]� �U�@D��tR��^]� V��^]� �����������̡�@@�@0�����U��V�u���t�Q�@@�@�Ѓ��    ^]����������U��V�@@��@V�ЋЋE����t��#��СR�@@V�@�Ѓ�^]� �U���u �E������   �$�u���   �u�u�u��]� ����������U�����   ���   ]����������̡Q�@H���   �Ѓ�������������U���u�@HQ��d  �Ѓ�]� �̡�@@�@T�����U���@@�@X]�����������������U���@@�@\]����������������̡�@@�@`�����U���@@�@d]�����������������U���@@�@h]�����������������U���@@�@l]�����������������U���@@���   ]�������������̡�@@�@t����̡�@@�@x�����U���@@�@|]����������������̡�@@���   ��U���@@���   ]�������������̡�@@���   �����   �@t��U���@@���   ]��������������U���@@���   ]��������������U���@@���   ]��������������U���@@���   ]��������������U���@@���   ]��������������U���@@���   ]��������������U���@@���   ]��������������U��V�u���t�Q�@@�@�Ѓ��    ^]���������̡�@@�@0�����U��j�@@�M�@4Qj �Ѓ�]����U��j�@@�M�@4Qh   @�Ѓ�]�U���u�@@�u�@4j �Ѓ�]���̡�@|� ������U��V�u���t�Q�@|�@�Ѓ��    ^]���������̡�@|�@ �����U��V�u���t�Q�@|�@(�Ѓ��    ^]����������U���@ �@H]�����������������U��}qF uGW�}��t>��u���   �ϋ@D�С�u�@@�@,�Ћ���ЋAW�u�@p����_]������������U���@��T  ]��������������U��S�@@V�@,W�u�Ћ�u�I@�؋I,�ы���yh��hE  �ˋ�����Ph��hE  �����P��T  �Ѓ�_^[]�����̡Q�@D�@$�Ѓ����������������U��j �@D�u� �Ѓ�]��������U��V�@@�u�@�6�Ѓ��    ^]��������������̡Q�@D�@�Ѓ���������������̡Q�@D�@�Ѓ���������������̡Q�@D�@(�Ѓ���������������̡Q�@D�@�Ѓ����������������U���@D� ]��U��V�@@�u�@�6�Ѓ��    ^]��������������̡Q�@D�@(�Ѓ���������������̡Q�@D�@�Ѓ���������������̡Q�@D�@(�Ѓ���������������̡Q�@D�@�Ѓ����������������U���u�@Dh2  � �Ѓ�]�����U��V�@@�u�@�6�Ѓ��    ^]��������������̡Q�@D�@(�Ѓ���������������̡Q�@D�@�Ѓ���������������̡Q�@D�@(�Ѓ���������������̡Q�@D�@�Ѓ���������������̡Q�@D�@(�Ѓ���������������̡Q�@D�@�Ѓ���������������̡Q�@D�@�Ѓ����������������U��j �@D�u� �Ѓ�]��������U��V�@@�u�@�6�Ѓ��    ^]��������������̡Q�@D�@(�Ѓ���������������̡Q�@D�@�Ѓ����������������U���u�@Dh'  � �Ѓ�]�����U��V�@@�u�@�6�Ѓ��    ^]��������������̡Q�@D�@(�Ѓ���������������̡Q�@D�@�Ѓ����������������U���u�@DhO  � �Ѓ�]�����U��V�@@�u�@�6�Ѓ��    ^]���������������U�����@XQ� �M�Q�ЋM�~ f��~@f�A�~@��f�A����]� ���������������U�����@XQ�@�M�Q�ЋM�~ f��~@f�A�~@��f�A����]� ��������������U�����@XQ�@�M�Q�ЋM�~ f��~@f�A�~@��f�A����]� ��������������U����`�@XV�@WQ�M�Q�Ћ��E���   ���_^��]� �������������U���u�@XQ�@�Ѓ�]� �����U���u�@XQ�@�Ѓ�]� �����U���u�@XQ�@�Ѓ�]� �����U���u�@XQ�@�Ѓ�]� �����U���u�@XQ�@$�Ѓ�]� �����U���u�@XQ�@ �Ѓ�]� ����̡j �@Dh�  � �Ѓ�����������U��V�@@�u�@�6�Ѓ��    ^]��������������̡Q�@D�@(�Ѓ���������������̡Q�@D�@�Ѓ����������������U���u�@D�u�@Q�Ѓ�]� �̡j �@Dh:  � �Ѓ�����������U��V�@@�u�@�6�Ѓ��    ^]���������������U�����E�    �E�    ���   �U��@Rj�����#E���]�����������̡j �@Dh�F � �Ѓ�����������U��V�@@�u�@�6�Ѓ��    ^]���������������U��E����u��]� �E���E�    ���   �U��@Rj������؋�]� ̡j �@Dh�_ � �Ѓ�����������U��V�@@�u�@�6�Ѓ��    ^]����������������    �A    �A    �A    �����V��V�G���FP�>�����F    �F    ^������������U��S�]V��W�~�    �    �F    �F    �CV;C��   ����W�����F    �F    �hg�@jI���   j�Ѓ������   �hg�@jN���   j�Ѓ����uV�������_^[]� ��F   �F   ����C�A��C�A�_�    ��^[]� �>��W�8���F    �F    �hg�@jI���   j�Ѓ����tZ�hg�@jN���   j�Ѓ�����X�����F   �F   ����C�A��C�A��C�A��    _��^[]� �����U��V�u���    �F    �F    �F    �  ��^]� U��V�u���  ��^]� �����������U��SV��V�C���FP�:���]���F    �F    ��t(�hg�H��    jIP���   �Ѓ����u^3�[]� W�}��t;�hg�H��    jNP���   �Ѓ��F��uV�����3�_^[]� �~_�^^�   []� �������������V��V����FP�~�����F    �F    ^������������U��SV��WV�R���^S�I���}���F    �F    ����   �? ��   �W����   �hg�H��    jlP���  �Ѓ����t<� t?�W��t8�hg�H��    jqP���  �Ѓ����u���%���_^3�[]� �G�F�G�F��P�7�6�+  �����t�F��P�wQ�z+  ��_^�   []� �����������U��SV��WV�R���~W�I�����} �F    �F    ��   �]����   �hg�@��    ���  h�   Q�Ѓ����t?�} tJ�U��tC�hg�H��    h�   P���  �Ѓ����u���)���_^3�[]� �E�F�,�F   �hg�@h�   ���  j�Ѓ����t���    P�u�^�6�g*  �M����t�F��PQ�7�N*  ���   _^[]� ��_^�   []� ����������������    �A    �A    �A    �����U������   �U��V�HWW�3��<��D$�|$@�L$}
��_^��]� ����  �0�U�f(ύ@�F�~ʍ@f(��D��,��t��\D��D$�\t��8�L$(�|$ �T$�\$0�\��D$8����   ��������f(ƍ@f(��$��T��\T��\��\��\\����Y��Y��Y��Y��\�f(��Y��Y��XL$(�\�f��\$0�\��L$(�Xl$�Xt$ �l$f�f(��D$ f�O�f����T$W��(��YL$(�YD$ �}f�?�X�f(��Y�f�f��X��@6  �T$(�\$ f(�W�f.͟��Dz�L$f(�f(�f(��&��b�^��L$f(�f(��Y��Y��Y�f�gH�%cfT�fT�f/�f�wPf�GX��   f(�fT�f/���   �GH�WX�gP(��Y�(��Y��\��Y��\�f�_�\�f�O f�g(�OX�P�Y(�W�gH(��YG (��YWP�\�(��YG(�Yg �Y�f�0�\��\�f�_8f�g@�)  �WPfT�f/��_X��   �OH�Y�f(��Y��\��\��Y�f�Gf�_ �\�f�O(�(�G �YGX�YP�O�wH(��Y_X�YOP�\�f(��YG(�Yw f�0�\��\�f�_8f�w@�   f(��Y�(��Y��\��GH�Y�f�O0�\��\�f�_8f�G@�oP�X�Y8�OH�w0(��YG@(��Y_@�YO8�\�(��YGX�Y�f��\��\�f�_ f�w(�D$`WP�����U���D$�   ���W�3�3Ʌ�~w��r]�p��W�W�%  �yH���@��+���    �o���f���oD��f��;�|�f��fo�fs�f��fo�fs�f��f~ϋt$;�}�F<�A;�|���t$�M��u�A0�D$(���q �@�D$    ���d��\��Y�f(��YI�D$(�Y��X	�D��Xq�@�X��AH�Y��X��A8�Y��L$ �I(�X��AP�Y��Y��T��X��A@�XI�Y��$��X��AX�Y�(��YY�X�(��YA0�Xf�L$X�L��D$�X�(��YAH�@���X�(��YA8�YQ@�\$(��YY �Ya(�D$�XY�Xa�X�(��YAP�YIX�X��X��X��\$0f�d$8���  3�������|$�D$(׋��@�,��T��L�f(��Ya(��YA0�X!f(��YY �Yi(�X��XY(��YAH�Xi�D$@�X�(��YA8�YQ@�D$�X�(��YAP�YIX�X��T$0�X�(��X�f(��\��\��\�f�\$0�YL$�YD$ �Y��X��~D$�D$ �~D$8f�D$X�X�f�f�d$f�l$8�X�;D$������|$@�D$@_^��]� ������������U�������������U�   @t������@��wg�$��o�E� ����E� ���]� �
�E��E�J�]� �J�E��E�J�]� �J�E��E�J�]� �J�E��E�
�]� ��Roho{o�o�o����U��S��V�����%���W��   @t�����ʃ��};�t�����t�u�����t��u;�t?�����t7�΁����Eǃ��t����   �_�^�[]� ��   ���Ё�   @�_^[]� �U�������AW�SVf(�f(�f(�W�L$�\$�T$ �D$���L  �9�u������Ш�)  ���������U��Z�@�[�<��l��\<��\l�;Zuc�\��B�\\��@�d��\d��T��\T��4��\4�f(��Y�f(��Y��Y��\�f(��Y��\��Xd$(��d�d��B�\d��@�B�@�T��\��\\��\T��4��\4�f(�f(��Y��Y��Y��\�f(��Y��\��X\$�XL$�Y��Y��\$�L$�\��Xt$ (��T$ ���L$�����f(��Y�f(��Y��X�f(��Y��X���-  f(�W�f.П��D�Ez� �@�@_^[��]� ��b�^�_^[(��YD$� (��YD$�@�D$�Y��@��]� ���������U���<�`g�5hg�A3�f�f�f�f��E��M��}��u��m��e�U�E����  S�V�uW�������Ш�v  ���������M��@��tn��f/�v	f(��E��\�f/�v	f(��M��\�f/�v	f(��}�f/�v	f(��u��T�f/�v	f(��m�f/�vIf(��>�~4��~l��~d�f�f�f�   �u��m��E��M��}ԉU��e�A�@��tn��f/�v	f(��E��\�f/�v	f(��M��\�f/�v	f(��}�f/�v	f(��u��T�f/�v	f(��m�f/�vIf(��>�~4��~l��~d�f�f�f�   �u��m��E��M��}ԉU��e�y���tn��f/�v	f(��E��\�f/�v	f(��M��\�f/�v	f(��}�f/�v	f(��u��T�f/�v	f(��m�f/�vIf(��>�~4��~l��~d�f�f�f�   �u��m��E��M��}ԉU��e�A;�t0�@�Mč�P�  �U��e��m��u��}��M��Eă��M��m���_^[��tb�Ef(��X�f(��X��Xgf(��X��Y��Y��Y�f�f�Pf�H�\0�\h�\`�Ef�0f�hf�`��]� �EW�f� f�@f�@�Ef� f�@f�@��]� ��������̋Q3���|�	��t��~�    t@��Ju��3�����������U��QV�u��;�}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}���x(���t"�v3Ʌ�~�I ���%���;�tA��;�|�_���^]� _��^]� ���������U��SV�q2ۅ�~:�W�}�
����%���;�u��   @u�����t	�   ���3�
؃�Nu�_��^��[]� �������������V�q3҅�~�	�d$ ��   @u	�����tB��Nu��^�����V�q3҅�~�	�d$ ����ШtB��Nu��^�����������U���V��3�9N~�A�d�����;N|��N��~jS�   3�W�U��]�����x9���������;�}*������<����������;�u��   ��@;F|ۋU��]��NB���B��]��U�;�|�_[^��]�����������h$jh_� �  ����uË@����U��V�u�> t/h$jh_� �  ����t��M�@�MQ�Ѓ��    ^]���U��Vh$jh_� ���Y  ����t�@��t�u����^]� 3�^]� ��������U��Vh$jh_� ���  ����t�@��t�u����^]� 3�^]� ��������U��Vh$jh_� ����
  ����t�@��t�u���u�u��^]� 3�^]� ��U��Vh$jh_� ���
  ����t�@��t�u����^]� 3�^]� ��������U��Vh$j h_� ���Y
  ����t�@ ��t�u����^]� 3�^]� ��������U��Vh$j$h_� ���
  ����t�@$��t�u����^]� 2�^]� ��������Vh$j(h_� ����	  ����t�@(��t��^��3�^������Vh$j,h_� ���	  ����t�@,��t��^��3�^������U��Vh$j0h_� ���y	  ����t�@0��t�u����^]� 3�^]� ��������U��Vh$j4h_� ���9	  ����t�@4��t�u���u��^]� ���^]� ����Vh$j8h_� ����  ����t�@8��t��^��3�^������U��Vh$j<h_� ����  ����t�@<��t�u����^]� ���������������U��Vh$j@h_� ���  ����t�@@��t�u����^]� ���������������U��Vh$jDh_� ���I  ����t�@D��t�u����^]� 3�^]� ��������U��Vh$jHh_� ���	  ����t�@H��t�u����^]� ���������������Vh$jLh_� ����  ����t�@L��t��^��3�^������Vh$jPh_� ���  ����t�@P��t��^��3�^������Vh$jTh_� ���l  ����t�@T��t��^��^��������Vh$jXh_� ���<  ����t�@X��t��^��^��������Vh$j\h_� ���  ����t�@\��t��^��^��������U��Vh$j`h_� ����  ����t�@`��t�u���u��^]� 3�^]� �����U��Vh$jdh_� ���  ����t�@d��t�u���u��^]� 3�^]� �����U��Vh$jhh_� ���Y  ����t�@h��t�u���u�u�u�u��^]� ���U��Vh$jlh_� ���  ����t�@l��t�u���u�u��^]� 3�^]� ��U��Vh$jph_� ����  ����t�@p��t�u���u��^]� 3�^]� �����U��Vh$jth_� ���  ����t�@t��t�u���u��^]� 3�^]� �����U��Vh$jxh_� ���Y  ����t�@x��t�u���u��^]� 3�^]� �����U��Vh$j|h_� ���  ����t�@|��t�u����^]� 3�^]� ��������U��Vh$h�   h_� ����  ����t���   ��t�u���u��^]� 3�^]� ���������������U��Vh$h�   h_� ���  ����t%���   ��t�u���u�u�u�u�u��^]� ���^]� ��U��Vh$h�   h_� ���6  ����t%���   ��t�u���u�u�u�u�u��^]� ���^]� ��U��Vh$h�   h_� ����  ����t���   ��t�u���u�u�u��^]� 3�^]� ���������U��Vh$h�   h_� ���  ����t���   ��t�u����^]� 3�^]� ��U��Vh$h�   h_� ���V  ����t���   ��t�u����^]� ���������U��Vh$h�   h_� ���  ����t���   ��t�u���u��^]� 3�^]� ���������������U��Vh$h�   h_� ����  ����t���   ��t�u���u�u��^]� 3�^]� ������������U����M�U�E�R�X�A�\B�\��\Y�Y �Y�Y�X��X��U��E���]�����U��h$�uh_� �+  ��]�������U��y0 �Etr��f/�v�	�H�Af/�v�I�H�Af/�v�I� f/Av�A�@f/A v�A �@f/A(vJ�A(]� �~ f�A�~@f�A �~@f�A(�~Af��~A f�A�~A(f�A�A0   ]� �������������U��Q���   �@X�Ћȃ���u]� ��u�@|�u�@Q�Ѓ�]� ����U��Q���   �@X�Ћȃ���u]� ��u�@|�u�@8Q�Ѓ�]� ����U��UV��j ��j �@j �@R�Ѓ��F��^]� ���̡V�@j �@j ��j �6�Ѓ��F^�U��V��N��u3�^]� �Q�u�@�u�@�6�Ѓ��F�   ^]� ������U��M�EQ��Ej�u�A�d����]���������������̸   �����������U��V�u��t���u6j�u�e������u3�^]Ë������ȅ�t��t��E3�;AOʋ�^]�������U��EHV����   �$�D��   ^]á4@�4����   �u蔓����=�6  }�����^]Ëu��t�hpgjmh<j��������tl���ʓ���0��tfV���Y����   ^]��u�u�����������H^]�^]�!����4u.�d����/s���50��t���^���V�x������0    �   ^]Ã��^]Ðp�����h�=�߄����U���Mu�E�(�E�,�   ]� ���������������U��h8jh�f �\�������t
�@��t]�����]�������U��Vh8jh�f �+���������t=�~ t7�u8�E�u4�u0�u,�u(����P�?����u�F�Ѓ�4�M���j�����^]ÍM����Z�����^]������U��h8jh�f ��������t
�@��t]��3�]��������U��h8jh�f ��������t
�@��t]��3�]��������U��h8�uh�f �[�����]������̃��\$�D$%�  =�  ��  �<$f�$f��f����  f$f�f(�fT�gf/�h�p  �8  f/�hsgf/�h��  f(�fY�f(�fY�f(-�hfY�fX-�hfY�fX-�hfY�fX-ph�Y�f(�f���X��Y��\Ń��f/�h��   f(�fY�f(�fY�f(-`hfY�fX-PhfY�fX-@hfY�fX-0hfY�fX- hfY�fX-hfY�fX- hfY�fX-�g�Y�f(�f���X��Y��\Ń���~�fW�f/�hsO�~�h�~-�h�~��X�fs�,f��f~؍@�~,Ũ��~��\��Y��X�h�^�f���   �~��~�h�^�f��~Ř��~$Š�f(�fY�f(�fY�f(-�hfY�fX-�hfY�fX-�hfY�fX-ph�Y�f(�f���X��Y��\��\��\�fVƃ��f/�hu	f$���f/ isf$�Y҃��f$f�g�Y҃���~��~�gfT�f.�z�D$��fi�X��g��ú�  ���T$�ԃ��T$�T$�$��  fD$���f�$�&  �$�~$��ÍI �������̃��\$�D$%�  =�  u�<$f�$f��f���d$�n  f��f%�f-00f=��6  fPq�Y�fXq�-��X�fpq�\�f(`q�Y�fɁ�v ����?f(-@q�i���fY��\��Yxq�\�fxf����\�fY�f\�f(5 q�Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-0q�Y fX5qfY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X��X�f(��f��f%�f��f�q�\�f(�Ã�f�$�  �$�~$����������̃��\$�D$%�  =�  u�<$f�$f��f���d$�{  f��f%�f-00f=��6  f z�Y�fz�-��X�f z�\�f(z�Y�fɁ� v ����?f(-�y��q���fY��\��Y(z�\�fxf����\�fY�f\�f(5�y�Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-�y�Y fX5�yfY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X��X�f(��,f��f=�u	�Y@z�f0z�Y��\��Y8zÃ�f�$��  �$�~$��ÍI Q�dz��  Y�U��V��������EtV�3���Y��^]� U���   �} t�I(  ��]øE�� �%�����������f��̴� 6��$��jh���H<  �E��uz�0  ��u3��F  �",  ��u�0  ����;  �`��1�97  �H�0  ��y�e,  ���w3  ��x �5  ��xj ��-  Y��u�D��   ��2  �Ʌ�ue�D��~�H�D�e� �=� u�-  �n,  �u��u��2  ��+  �0  �E������   �   �u��u�=(�t��+  ��p��u^�5(�C7  Y��u[h�  j�:  YY���������V�5(�97  YY��tj V�Z*  YY�`��N��V�t  Y�������uj �u)  Y3�@�*;  � U��}u�h5  �u�u�u�   ��]� jh���:  3�@�u��u95D��   �e� ��t��u5�lz��t�uV�u�щE����   �uV�u�����E����   �]SV�u�m������}��u(��u$SP�u�U���SW�u������lz��tSW�u�Ѕ�t��u*SV�u�������#��}�t�lz��tSV�u�Ћ��}��E��������&�M�Q�0�u�u�u�   ��Ëe��E�����3���9  �U��}u�uj �u�G����u�u��&  YY]�U��} t-�uj �5��`��uV�;  ���`P�;  Y�^]�U��V�u���woSW����u��  j�>  h�   ��)  ��YY��t���3�AQj P�`����u&j[9�tV�q;  Y��u���;  ��
;  ���_[�V�P;  Y��:  �    3�^]��̋T$�L$��t�D$�%�s�L$W�|$��]�T$���   |�%��.;  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�;� u����=  �WV�t$�L$�|$�����;�v;��h  �%�s��  ���   ��  ��3Ʃ   u�%���  �%� ��  ��   ��  ��   ��  ��s����v����s�~���vf����   tc����   foN�v�fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�   foN��v��I fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�VfoN��v���fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v��|�o���vf�����s����v����s�~���vf����X�����   u������r*��$�X���Ǻ   ��r����$�l��$�h���$���|���̔#ъ��F�G�F���G������r���$�X��I #ъ��F���G������r���$�X��#ъ���������r���$�X��I O�<�4�,�$�����D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�X���h�p�|����D$^_Ð���D$^_Ð���F�G�D$^_ÍI ���F�G�F�G�D$^_Ð�t1��|9���   u$������r����$��������$����I �Ǻ   ��r��+��$����$�����,�T��F#шG��������r�����$����I �F#шG�F���G������r�����$�����F#шG�F�G�F���G�������V�������$����I ��������ȖЖؖ��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��������0��D$^_Ð�F�G�D$^_ÍI �F�G�F�G�D$^_Ð�F�G�F�G�F�G�D$^_Í�$    W�ƃ�����   �у���te��$    �fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tO������t��    fof�v�Ju��t*����t���v�Iu�ȃ�t��FGIu���    X^_Í�$    ���̺   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y�����Vjj �0  YY��V� `��1��1��ujX^Ã& 3�^�jh���1  ��$  �e� �u�#   Y���u��E������   ���1  Ëu��$  �U��QSV�5`W�5�1���5�1�E��֋؋E�;���   ��+��O��rvP��7  ���GY;�sG�   ;�s�Ƌ]��;�rPS�{0  YY��u�F;�r>PS�g0  YY��t1��P��� `��1�u� `�KQ�� `��1�E�3�_^[��U���u����������YH]���WV�t$�L$�|$�����;�v;��h  �%�s��  ���   ��  ��3Ʃ   u�%���  �%� ��  ��   ��  ��   ��  ��s����v����s�~���vf����   tc����   foN�v�fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�   foN��v��I fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�VfoN��v���fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v��|�o���vf�����s����v����s�~���vf����؜����   u������r*��$�؜��Ǻ   ��r����$���$����$�l����(�L�#ъ��F�G�F���G������r���$�؜�I #ъ��F���G������r���$�؜�#ъ���������r���$�؜�I Ϝ���������������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�؜��������D$^_Ð���D$^_Ð���F�G�D$^_ÍI ���F�G�F�G�D$^_Ð�t1��|9���   u$������r����$�t������$�$��I �Ǻ   ��r��+��$�x��$�t������ԝ�F#шG��������r�����$�t��I �F#шG�F���G������r�����$�t���F#шG�F�G�F���G�������V�������$�t��I (�0�8�@�H�P�X�k��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�t������������D$^_Ð�F�G�D$^_ÍI �F�G�F�G�D$^_Ð�F�G�F�G�F�G�D$^_Í�$    W�ƃ�����   �у���te��$    �fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tO������t��    fof�v�Ju��t*����t���v�Iu�ȃ�t��FGIu���    X^_Í�$    ���̺   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y����������������̃��\$�D$%�  =�  ��   �<$�$������   f����%�  =�  t0��% �  u�Q����f�$�<$ uP�� �  uHf���� u>�ً���u$f��%��  uf��%��  uf�� %��  t�f�$�L$��  ��$    �D$  ���1   ���T$�ԃ��T$�T$�$�  fD$���f�$�R0  �$�~$��Ë�j�4  Y��tj�4  Y��u�=Puh�   �1   h�   �'   YY�U��M3�;���t
@��r�3�]Ë���]�U����  �� 3ŉE�V�uWV������Y���y  Sj�4  Y���  j�4  Y��u�=P��   ���   �A  h�h  hX�2  ��3ۅ��/  h  h�Sf���$`��  ��uh@�Vh��i2  ������   h��2  @Y��<v5h��2  �E��-�j��hp�+�VQ�2  ������   hx�h  �XV�1  ������   Wh  V�1  ����u{h  h��V�H3  ���Wj��`����tI���tD3ۋˊO�����f9Ot	A���  r�S�����P�����P�]��0  YP�����PV� `[�M�_3�^������SSSSS�>0  ��4  ��tj��4  Y�� t!j腵  ��tjY�)jh  @j�.  ��j�  �U��E��]�U���(3��E��E�9�t�5�1�`����&��E��   V;���  ��  ���  ��   jZ+���   H��   ����   H��   ����   HtN��	�#  �E�   �E�H��E�u� �E�]�� �E��]�P��]���Y����  �O(  � "   ��  �E�D��E�u� �E�]��E�   � �E��]�P��]���Y�  �E�   �E�D���E�<��V  �U��E�<��l����E�8��;  �U��E�8��Q����E�H�놃�tfHtWHtHHt/���  ��	t���8  �E�L���   �E�T���   �E�H��E�u� ���   �E�H���   �E�   �������E���   �E�   �E�\������������   �$���E�8���E�<���E�D���E�d���E�l��u����E�t��i����E�|��]����E܄��E�u� �M��� �E�]�� �]��.�E܈����E܌����Eܐ��E�u� �E�]�� �]���E��]�P�E�   ��Y��u�q&  � !   �E��^�Ë�E�N�W�`�i�u�����פˤ������¥�= 1 ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU��4  ��= 1 t2���\$�D$%�  =�  u�<$f�$f��f���d$u�4  ���$��9  �   ��ÍT$�m9  R��<$t6f�<$t�-������=@ ��9  �   �� �9  �9  �&��� u�|$ u����-���   �t���뻸   �=@ �V9  �   �� �O:  Z������̃= 1 ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU�i:  ��= 1 t2���\$�D$%�  =�  u�<$f�$f��f���d$u�:  ���$�8  �   ��ÍT$�M8  R��<$tPf�<$t�-��������z�=@ �|8  �   �� �y8  �-����������z���������7  ���� u�|$ u����-���   �=@ �'8  �   �� � 9  Z�������̃= 1 ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU��:  ��= 1 t2���\$�D$%�  =�  u�<$f�$f��f���d$u�:  ���$�r7  �   ��ÍT$�7  R��<$tPf�<$t�-��������z�=@ �L7  �   �� �I7  �-����������z��������6  ���� u�|$ u����-���   �=@ ��6  �   �� ��7  Z�������̋T$�L$��   u@�:u2��t&:au)��t��:Au��t:au������uҋ�3���������Ë���   t���:u����t���   t�f���:u΄�t�:auń�t����jh���  j�^;  Y�e� �u�F��t0�����M��t9u,�A�BQ�$���Y�v����Y�f �E������
   ��  Ë���j�f<  Y�U��V��M�F ��uf�*  �ЉV�Jl��Jh�N�;�
t���Bpu�@  ��F;@t�N���Apu�~C  �F�N�Ap�u���Ap�F�
���A�F��^]� U��j �u�u�u�u�u�u�   ��]�U��E��et_��EtZ��fu�u �u�u�u�u��  ��]Ã�at��At�u �u�u�u�u�u�s  �0�u �u�u�u�u�u�   ��u �u�u�u�u�u��  ��]�U���,SVWj0X�u�ȉM��M��E��  3������}��y���u��t�M��u	�<   j��G�;�w�*   j"_�8��&  ��  �U��Z�E����%�  =�  uy3�;�uu���;�t�A�j WP�^SR�  ������t� �  �;-u�-F�}j0X�������$�x�F�FjeP�H  YY��t�����ɀ����p��@ 3��O  3���   ��t�-F�} �]j0X�����$�x��ۈF�J�����'��  �3���]�u'j0X�F�B�
%�� ���u3��E���E��  ��F1����F�M��u� ��Eԋ��   � � ��B%�� �E�w	�: ��   �e �E��   �M��~S��R#E#ыM��Ɂ��� �YL  j0Yf�����9vËM�U��E���E�E�����FO�M�E�f��y�f��xW��R#E#ыM��Ɂ��� �L  f��v6j0�F�[���ft��Fu�H��]�;E�t���9u��:��	�����@���~Wj0XPV�&�������E�8 u���} �U����$�p���R�4�K  ��3��ځ��  #�+M��x;�r	�F+����F-������ۋ��0;�|A��  ;�rPRSQ�[J  0�F3��U�;�u;�|��drPjdSQ�8J  0�F�U�3�;�u;�|��
rPj
SQ�J  0��U�F�]�3���0��F���}� t�M܃ap���_^[��U��j �u�u�u�u�u�T  ��]�U����M�SW�u �F����]��t�} w	��  j��U3����ǃ�	9Ew��  j"_�8�#  ��   �} t �M3�����P3��9-���P��  �UYY�EV�8-��u�-�s��~�F��E�F���   � � �3�8E�������9Et��+�Eh��PV�;5  ����ut�N9}t�E�U�B�80t-�RJy���F-jd[;�|��� Fj
[;�|��� F V�� ^t�90uj�APQ�������}� t�M��ap���_[��WWWWW�"  �U���,�� 3ŉE��ES�]VW�}j^V�M�Q�M�Q�p�0�G  ����u�x  �0�="  ���t�u��u
�a  j^����;�t3��}�-����+�3�����+ȍE�P�CPQ3Ƀ}�-��3�������P�D  ����t� ��u�E�j P�uSVW��������M�_^3�[������U����ES�@V�uH�M�E��!����u��t�} w�  j[��}!  �   3�W�}8]t�M�;�u�U3��:-���f�00 �E�8-u�-F�@��jV�  Y�0YF����~JjV�  �E�Y���   Y� � ��EF�@��y&8]t�������;�|��WV�`  Wj0V�.�����_�}� t�M�ap�^��[��U���,�� 3ŉE��ESW�}j[S�M�Q�M�Q�p�0��E  ����u��  ��   ���lV�u��u�  ��s   ���S���;�t3��}�-����+ȋ]�E�P�E��P3��}�-Q���P�C  ����t� ��u�E�j PSVW�i�����^�M�_3�[�������U���0�� 3ŉE��ESW�}j[S�M�Q�M�Q�p�0�?E  ����u�  ���  ���   V�u��u��  ��  ���   �E�H3Ƀ}�-�E�������9;�t��+��M�Q�uPS�PB  ����t� �S�E�H9E������|+;E}&��t
�C��u��C��u�E�jP�uVW��������u�E�jP�u�uVW�Q�����^�M�_3�[�������U��j �u�   YY]�U���W�u�M��u����U�}��
��t���   � � :�tB�
��u��B��t4�	<et<EtB���u�V��J�:0t����   ��:uJ�BF���u�^�}� _t�E��`p���U��j �u�u�u�   ��]�U��QQ�} �u�ut�E�P��A  �M�E���E��A��EP�DB  �M�E�����U��j �u�   YY]�U����M�V�u�����u�P�b?  ��e�F�P��=  ��Yu��P�E?  Y��xu���E�����   � � �F���ȊF��u�^8E�t�E��`p���U��E�������Az3�@]�3�]�U��W�}��tV�uV�  @P�>VP�������^_]�Vh   h   3�V�KD  ����u^�VVVVV�N  �V3��� � `�� ����(r�^�U��V��  �����E  �V\W�}��99t�����   ;�r�   ;�s99t3Ʌ��  �Q���  ��u�a 3�@��   ��u�����   �ES�^`�F`�y��   j$_�F\���d� ���   |�9�  ��~du�Fd�   �   �9�  �u	�Fd�   �u�9�  �u	�Fd�   �d�9�  �u	�Fd�   �S�9�  �u	�Fd�   �B�9�  �u	�Fd�   �1�9�  �u	�Fd�   � �9� �u	�Fd�   ��9� �u�Fd�   �vdj��Y�~d�	�q�a ��Y�^`���[�3�_^]�U��csm�9Eu�uP����YY]�3�]�jh0��  �u���   �~$ t	�v$�����Y�~, t	�v,�����Y�~4 t	�v4�����Y�~< t	�v<�����Y�~@ t	�v@�����Y�~D t	�vD����Y�~H t	�vH����Y�~\��t	�v\����Yj�-  Y�e� �~h��tW�4`��u��@tW�f���Y�E������W   j�[-  Y�E�   �~l��t#W�2  Y;=�
t���
t�? uW�0  Y�E������   V����Y��  � �uj�h.  YËuj�\.  Y�U��(���t'V�u��uP�T  ��(Yj P�c  YYV����^]�V�   ����uj�  Y��^�VW�`�5(���  ��Y��uGh�  j��  ��YY��t3V�5(�  YY��tj V�%   YY�`�N���	V�?���Y3�W�,`_��^�jhX��  �u�F\���f 3�G�~�~pjCXf���   f���  �Fh@���   j��+  Y�e� �vh�0`�E������>   j��+  Y�}��E�Fl��u��
�Fl�vl�.  Y�E������   �g  �3�G�uj��,  Y�j��,  Y��  �,  ��u�c   3��h���  Y�(���t�Vh�  j�  ��YY��t-V�5(��  YY��tj V�����YY�`�N��3�@^��   3�^á(���tP�Z  �(�Y�'+  U��Q�E�PhP�j �<`��thh��u��@`��t�u����U���u�����Y�u�8`�VW�5�1�`�5�����t�> t�6�|���Y��u�5�SV�i����5�3�Y����t9t�6�K���Y��u�5�V�9����5����(����5��������������t9�1tW�����Yj�� `��1�� ��tP�����Y�� �� ��tP�����Y�� �5@�4`[��u�@�@;�tP����Y�5@_^�U��������u����Yh�   �   �jj j �1  ���U��=hz thhz�>  Y��t
�u�hzY����h(aha��   YY��uPVWh������Y�a�a����t�Ѓ�;�r�=�1 _^th�1�'>  Y��tj jj ��13�]�U��j j�u�   ��]�Vj � `��V��  V��  V�<���V�?  V�  V��>  ��^�	  U��V�u����t�Ѓ�;ur�^]�U��V�u3����u���t�у�;ur�^]�j�N(  Y�j�)  Y�jh���  j�0(  Y�e� �=���   ��   �E���} ��   �5�1�5`�֋؉]ԅ�tt�5�1�֋��]�}��}܃��}�;�rWj � `9t�;�rG�7�֋�j � `����5�1�5`�։E��5�1�֋M�9M�u9E�t��M�ى]ԉE����h<ah,a�����YYhDah@a�����YY�E������    �} u)��   j�(  Y�u�h����} tj�(  Y���  ��H`3Ʌ�������Ã%� �jdh���n  j��&  Y3ۉ]�j@j _W�5
  YY�ȉM܅�uj��E�Ph� �;(  ������U  ���=�1   ;�s1f�A 
�	��Y�a$��A$$�A$f�A%

�Y8�Y4��@�Mܡ��ƍE�P�X`f�}� �)  �E����  ��M���E���E�   ;�|�ȉM�3�F�u�9�1} j@W�v	  YY�ȉM܅���   ��1�M���}ԋE؋U�;���   �2���tX���tS� �tM�uV�L`�U���t8����������4���u܋��E؊ �Fh�  �FP�P`�F�U��M�G�}ԋE�@�E؃��U�놉��=�1���   ;�s$f�A 
�	��Y�a$�f�A%

�Y8�Y4��@�M���F�uЋM������]ԃ���   ����5��u܃>�t�>�t�F��F�   �F���uj�X�
�C�������P�`�����tE��tAW�L`��t6�>%�   ��u�F@���u	�F�Fh�  �FP�P`�F�"�F@�F������!��t
���@����C�<����E������   3��	  �j�%  Y�VW���>��t7��   ;�s"���� tW�T`���@��   �G�;�r��6� ����& Y�����|�_^�U��QQ�=�1 u�*  SVWh  ��3�WS���\`�5�1�=���t8u���E�P�E�PSSV�[   �]��������?sE�M����s=��;�r6R�*  ��Y��t)�E�P�E�P��PWV�   �E���H���=�3�����_^[��U��ES�]V�# �u�    �EW�}��t�8���E3ɉM�>"u3�����F�ȉM�"�5���t��G��E��PF�);  Y��t���t��GF�E��t�M��u�< t<	u���t�G� �N�e �> ��   �< t<	uF��> ��   �U��t�:���U�E� 3�B3��FA�>\t��>"u3��u�} t�F�8"u���3�3�9E���E���I��t�\G���u���tA9Mu< t8<	t4��t*��P�V:  Y��t��t��GF���G���tF��F�o�����t� G��-����U_^[��t�" �E� ]Ã=�1 u��'  V�5HW3���u����   <=tGV�N  FY����u�GjP��  ��YY�=���tʋ5HS�> t>V�  �>=Y�Xt"jS�  YY���t@VSP��   ����uH���> uȋ5HV�����%H �' ��1   3�Y[_^��5�������%� �����3�PPPPP�r  �U����� �e� �e� VW�N�@��  ��;�t��t	�У� �f�E�P�h`�E�3E�E��`1E��d`1E��E�P�``�M�3M�E�3M�3�;�u�O�@����u��G  ��ȉ� �щ� _^��U��QW�l`��3���tuV��f9t��f9u���f9u�SPPP+�P��FVWPP�t`�E���t7P�  ��Y��t*3�PP�u�SVWPP�t`��u	S�����Y3�W�p`���	W�p`3�[^_��U��@13� t�u��]�]�%�`U��D13� �ut��]���`]�U��H13� �ut��]���`]�U��L13� �u�ut��]���`]�U��QV�5p��y%��13�3� �u�tV�M�Q�Ѓ�zuF�5p3�����^��VWhx���`�5@`��h��W��3� h��W�@1��3� h��W�D1��3� h��W�H1��3� h��W�L1��3� hܞW�P1��3� h�W�T1��3� h�W�X1��3� h �W�\1��3� h4�W�`1��3� hT�W�d1��3� hl�W�h1��3� h��W�l1��3� h��W�p1��3� h��W�t1��3� �x1hȟW��3� h�W�|1��3� h�W��1��3� h$�W��1��3� h8�W��1��3� hT�W��1��3� hh�W��1��3� hx�W��1��3� h��W��1��3� h��W��1��3� h��W��1��3� hĠW��1��3� hؠW��1��3� h�W��1��3� _��1^�U���u��`P��`]�U��j �|`�u�x`]�U��VW3�j �u�u�5  ������u'9�vV��`���  ��;�v������uË�_^]�U��SVW�=�3��u�m�����Y��u%��t!V��`�=����  ��;�v������u�_^��[]�U��VW3��u�u�Q4  ��YY��u,9Et'9�vV��`���  ��;�v������u���_^]�VW����������t�Ѓ�;�r�_^�VW����������t�Ѓ�;�r�_^���h��d�5    �D$�l$�l$+�SVW�� 1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q��������U���S�]VW�{3=� �E� �E�   ��s���t�O�30�9����O�G�30�)����E�@f��   �E�E�E�E�C��C�E������   �@�@�L������E���t{���  ��M����~   ~h�E�8csm�u(�=$1 th$1�/  ����tj�u�$1���U�M��  �E�U�9Pth� V����  �E�X����tu�f�M��É]�����]�����tG�!�E�    ��{�t6h� V�˺�����  ����t�O�30� ����O�W�32�����E�_^[��]ËO�30������O�G�30������M��֋I�  ��������u��Ã��U��V������MQ��    Y���   �0^]�������u��Ã��U��M3�;ŀt'@��-r�A��wjX]Í�D���jY;��#���]Ëń]�U���5��`��t�u��Y��t3�@]�3�]�U��E��]Å�uf���fn�f`�fa�fp� SQ�ك���ux�ڃ���t0ffAfA fA0fA@fAPfA`fAp���   KuЅ�t7����t��I f�IKu���t����t
f~�IJu���t�AKu�X[��ۃ�+�R�Ӄ�t�AJu���t
f~�IKu�Z�^���U��%� ��S3�C	�j
�؊  ���  3ɋÉ��V�5�W�}�����_�O�W�E�   �5�t����   �5��E�   t����   �5�j3�X��u���^�N�V�E�   �5�t	���5�3�3���}���_�O�W�}�Genuu_�}�ineIuV�}�nteluM3�@3����_�O�W�E�%�?�=� t#=` t=p t=P t=` t=p u	���5�_^3�[��U���uj �u�u�u�   ��]�U��� �e� Wj3�Y�}��9Eu�>����    ��  ����x�EV�u��t��u�����    ��  ����S�����M�;�w�E��u�E��u�E�B   �u�u�P�u���0  ������t�M�x�E��  ��E�Pj �/  YY��^_��U����`j��.=  �u�6����= YYuj�=  Yh	 �����Y]�U���$  j諈  ��tjY�)���������5��=�f� f��f��f��f�%�f�-�����E ���E���E���������8  ������	 ���   ��   jXk� ǀ�   jXk� �� �L�jX�� �� �L�h���������U��} u�o����    �0  ���]��uj �5���`]���̃��$�]  �   ��ÍT$�  R��<$�D$tQf�<$t��  �   �u���=@ �3  �   � �0  �  �u,��� u%�|$ u���  �"��� u�|$ u�%   �t����-���   �=@ ��  �   � ��  Z�U���(  �� 3ŉE��}�Wt	�u��:  Y������ jL������j P�l�����������������0�����������������������������������������������f������f������f������f������f������f��������������E�������E������ǅ0���  �@��������E�������E�������E��������`��������P�1���Y��u��u�}�t	�u�
:  Y�M�3�_������U��E�]�U���5�`��t]���u�u�u�u�u�   �3�PPPPP��������j�b�  ��tjY�)Vj� �Vj�u���V������^ËL$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+��U��VW�}��t�M��t�U��u3�f��J���j^�0������_^]Ë�f�> t��Iu��t�+��f��Rf��tIu�3���u�f�����j"�U��V�u��t�U��t�M��u3�f������j^�0������^]�W��+��f��If��tJu�3�_��u�f�����j"��U��Ef���f��u�+E��H]�U��U�MV��u��u9Mu&3��3��t�E��t��u3�f���u��u3�f��K���j^�0������^]�SW�ً����u+��f�3�vf��t%Ou�� +��f��[f��tOtJu��u3�f���_[�{������u�E3�jPf�TA�X�3�f������j"�U��E��x!��~��u������]������    �`������]�U���$�� 3ŉE��ES� `VW�E�E3�W�E��Ӌ��u��i����E�9=��   h   Wh���`����u$�`��W�h  h���`�����S  h�V�@`���?  P��h(�V��@`P��h8�V��@`P��hL�V��@`P�ӣ ��thh�V�@`P�ӣ�u���`��t�E��tP��`9}�tjX�   9}�t�5�`j���`;�tO95 tGP���5 �E��ӋM�E��t/��t+�х�t�M�Qj�M�QjP�U��t�E�u�u��    �0�;�t$P�Ӆ�t�Ћ���t�;�tP�Ӆ�tW�Ћ��u�5�Ӆ�tV�u��u�W���3��M�_^3�[�V������5,�`�U��E�$�(�,�0]�j$h���O���3ۉ]�3��}؋u��Pt��jY+�t"+�t+�t^+�uH��������}؅�u����d  �E�$�$�^�w\V�S  YY���E� �V�ƃ�t6��t#Ht�����    �������E�,�,��E�(�(��E�0�03�C�]�P�`�E܃���   ��uj������tj ��  Y�e� ��t
��t��u�G`�EЃg` ��uA�Gd�E��Gd�   ��u/�H��щUԡL��;�}&��k��G\�d B�UԋH���j � `�M��E������   ��u �wdV�U�Y��u�]��}؅�tj �  Y�V�U�Y��t
��t��u�EЉG`��u�ẺGd3�������U��M�@�V�u9qt��k�E��;�r�k�U;�s	9qu���3�^]�U��E��t���8��  uP�ö��Y]�U��SVW3���   �;�+���jU�4����u�   ����ty�^���~;�~Ѓ�������_^[]�U��} t�u����Y��x=�   s	�ŀ�]�3�]�U�졬13� t3�QQQ�u�u�u�u�u�u��]��u�u�u�u�u�u����YP��`]�U��V�u3���t^�MSW�}jA[jZZ+��U�jZZ�f;�rf;�w�� ������f;�rf;Ew�� ����Nt
f��tf;�t�����_+�[^]�3��j
�~}  � 13����������U�������$�~<$�   ���~|$f�f(�fTP�f/x���  �U  f/h�snf/p���  f(�fY�f(�fY�f(- �fY�fX-�fY�fX- �fY�fX-���Y�f(�f���X��Y��\�f�|$�D$�f/`���   f(�fY�f(�fY�f(-��fY�fX-��fY�fX-��fY�fX-��fY�fX-��fY�fX-��fY�fX-��fY�fX-p��Y�f(�f���X��Y��\�f�|$�D$��~�fW�f/X�sO�~P��~-0��~��X�fs�,f��f~؍@�~,Ũ��~��\��Y��XH��^�f���   �~��~@��^�f��~Ř��~$Š�f(�fY�f(�fY�f(- �fY�fX-�fY�fX- �fY�fX-���Y�f(�f���X��Y��\��\��\�fV�f�D$�D$�f/8�u�D$�f/��s���������$�$���D$��������D$��~��~@�fT�f.�z�D$�������`�ú�  ���T$�ԃ��T$�T$�$�5������D$Ð���̀zuf��\���������?�f�?f��^���٭^�������剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�������剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp���������۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-����p��� ƅp���
��
�t�����������������������������ËT$��   ��f�T$�l$é   t�   �����   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   ��   Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t�{   Z��]   Z��,$Z����������������������   s��������������������������   v���������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�l+  ���E�f�}t�m���������������U�������$�~$�   ��fD$f��f%�f-00f=��B  fP��Y�fX��-��X�fp��\�f(`��Y�fɁ�v ����?f(-@������fY��\��Yx��\�fxf����\�fY�f\�f(5 ��Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-0��Y fX5�fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���+f��f%�f����f���\�fL$�D$����V����I ����U�������$�~$�   ��fD$f��f%�f-00f=��B  f ��Y�f��-��X�f ��\�f(��Y�fɁ� v ����?f(-��������fY��\��Y(��\�fxf����\�fY�f\�f(5���Y��\�fY�fY��\�f(�\�fX�X��\��Y�fY��Y�fY�fY�fX-���Y fX5��fY����XX�Y����X�fX�fh�\��\��XHfY��X��X��X��X��X�f��X΃��X�fd$�D$���I��f��f=�u�Y@�fD$�D$���f0��Y��\��Y8�fD$�D$��������U��V�u��t�U��t	�M��u������j^�0������^]�W��+���A��tJu�_��u�����j"��3���U��V�u�<�  uV�q   Y��uj�B���Y�4� ��`^]�VW� ��S���t�tS�T`S蠪���' Y����@|�[�> t�~u�6�T`����@|�_^�jh��������=� u葺��j����h�   ����YY�}�<�  u[j�����Y����u������    3��Aj
����Y�e� �<�  uh�  V�P`�4� �V����Y�E������	   3�@�����j
�7   Y�VW� �@�~u�>h�  �6���P`����@|�3�_@^�U��E�4� ��`]�����������SVW�T$�D$�L$URPQQh��d�5    �� 3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�R(  �   �C�d(  �d�    ��_^[ËL$�A   �   t3�D$�H3�� ���U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�'  3�3�3�3�3���U��SVWj Rhv�Q�>p  _^[]�U�l$RQ�t$������]� U��SV�50`W�}W�փx t�wx�֋��   ��tP�փ| t�w|�֋��   ��tP��jX�_�E�{�`	t�; t�3�֋E�{� t�{� t�s��֋E��H�Eu΋��   �   P��_^[]�U��SV�u3ۋ��   W��tf=8t_�Fx��tX9uT���   ��t9uP�W������   �&  YY�F|��t9uP�9������   �'  YY�vx�$������   ����YY���   ��tD9u@���   -�   P��������   ��   +�P�������   +�P�צ�����   �̦�������   =h	t9��   uP�'  ���   裦��YYjX���   �~�E��`	t���t�8 uP�x����3�q���YY�E�� t�G���t�8 uP�T���Y�E����H�Eu�V�>���Y_^[]�U��V�u����   SW�=4`V�׃~x t�vx�׋��   ��tP�׃~| t�v|�׋��   ��tP��jX�^�E�{�`	t�; t�3�׋E�{� t�{� t�s��׋E��H�Eu΋��   ���   Q��_[��^]�jh ���������������Npt"�~l t�����pl��uj �����Y���/����j�_���Y�e� �5�
�FlP�!   YY���u��E������   뼋u�j����Y�U��W�}��t;�E��t4V�0;�t(W�8�����Y��tV�����> Yu���
tV�O���Y��^�3�_]Ã=�1 uj��P  Y��1   3��U��E-�  t&��t��tHt3�]á��]á��]á��]á��]�U����M�j �w����E�%�  ���u��    ��`�,���u��    ��`����u�E���    �@�}� t�M��ap���U��S�]VWh  3��sWV�Ĥ��3��ȉ{�{��  ������{����@��+��  �7�FIu���  �   �9�AJu�_^[]�U���   �� 3ŉE�SV�uW������P�v��`3ۿ   ����   �È�����@;�r�����ƅ���� ��������Q���;�sƄ���� @;�v�����u�S�v������PW������PjS�*  S�v������WPW������PW��  S�.)  ��@������S�vWPW������Ph   ��  S�)  ��$����M�����t�L��������t�L ��������  ���  A;�r��Wj���  X+ˉ������������� ��w
�L�A �������w�L �A����������A��  ;�r��M�_^3�[�y�����jh ������S��������Opt�l t�wh��uj �W���Y�������j�����Y�e� �wh�u�;5@t6��tV�4`��u��@tV詡��Y�@�Gh�5@�u�V�0`�E������   뎋u�j�����Y�jh@��������������؉]��=����sh�u�����Y�E;F�n  h   �����Y�؅��[  ��   �E�ph���3��3S�u�G  YY���}���  �E��ph�4`���E�u�Hh��@t
Q�ܠ��Y�E�XhS�0`�E��@p��   ����   j����Y�u��C�� �C�� ��  �� �ΉM���}f�DKf�M� A��ΉM���  }�D��8A��u���   }��  ��@F���5@�4`��u�@=@tP����Y�@S�0`�E������   �1�}j�d���Y��#���u��@tS�����Y�����    �3��������U��� �� 3ŉE�SV�u�u�-�����Y�]���uV����Y3��  W3��ωM��9�H��   A��0�M�=�   r����  ��   ����  ��   ��P��`����   �E�PS��`����   h  �FWP�����^3�C����  9]�vO�}� �E�t!�P��t�����LA;�v����8 uߍF��   �@Iu��v��������  �^��~3��ȋ�����~����   9=� tV�����   ����   h  �FWP�H����U��k�0��X�E�8 ��t5�A��t+������   s��DD�AC;�v���9 u΋E�G���E��r��]�S�^�F   �W�������  j�N��L_f�f��R�IOu�V�<���Y3�_�M�^3�[�1�����U����u�M��˷���M��yt~�E�Pj�u�X%  ��������   �E�A���}� t�E��`p�����U��=! u�M�`�H��]�j �u����YY]�U����M�SW�u�N����]�   ;�s`�M�yt~�E�PjS��$  �M������   �X����t�}� ���   �t�E��`p�����   �}� t�M��ap����   �E�xt~-�����E�M���QP�i%  YY��t�Ej�E��]��E� Y��S���� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QW���   �E�P�"  ��$��u8E��{����E��`p��o�����u�}� �E�t%�M��ap���U��E���Ѐ}� t�M��ap���_[��U��=! u�M�A���w�� ��]�j �u����YY]��������U��W�=���   �}ww�U�����fn��p� ۹   #σ����+�3��of��ft�ft�f��#�uf��#���ǅ�EЃ������Sf��#���3�+�#�I#�[��ǅ�D�_���U��t93���   t�;�Dǅ�t G��   u�fn�f:cG�@�L�B�u�_�ø����#�f��ft �   #Ϻ������f��#�uf��ft@��f����t����뽋}3�������ك��E���8t3�����_��U��UV�uW�z��u�K���j^�0�������   �} v�M� ��~���3�@9Ew	����j"��S�^�0�Å�~���t��G�j0Z�@I���U�  ��x�?5|�� 0H�89t�� �>1u�B�S�����@PSV������3�[_^]�U���(�� 3ŉE�SV�uW�u�}�M������E�P3�SSSSV�E�P�E�P�-  �E�E�WP�"  �ȋE��(�u��t��uj�
�u��tj[�}� t�M��ap��M�_^��3�[�Ϛ����U���(�� 3ŉE�SV�uW�u�}�M��V����E�P3�SSSSV�E�P�E�P�
-  �E�E�WP�'  �ȋE��(�u��t��uj�
�u��tj[�}� t�M��ap��M�_^��3�[�C�����U��QQ�ES�PVW�x� �������  �� �  ����� �   ��}��E���t���  t�� <  �%��  �!��u��u�E!P!f�x�X��<  3����M���������]���E�s���x&�������������  �y�}�}��E�s�f�{_^[��U���0�� 3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���uЋ���f��,3  �u܉C�E��E��C�E�P�uV�o�����$��u�M�_�s^��3�[�������3�PPPPP�%�������������������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��U��M�E������#�V�u�����t$��tj j �<  YY�����j^�0��������Q�u��t	��;  ����;  YY3�^]�j����Y������������U��ES�H<�V�A�Y��3��W��t�}�p;�r	�H�;�r
B��(;�r�3�_^[]��������������U��j�h`�h��d�    P��SVW�� 1E�3�P�E�d�    �e��E�    h   �|   ����tT�E-   Ph   �R�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE� 3Ɂ8  �����Ëe��E�����3��M�d�    Y_^[��]�������U��E�MZ  f9t3�]ËH<�3��9PE  u�  f9Q��]�jh���S��������@x��t�e� ���3�@Ëe��E�����������h��� `�� �U��E�� ]á!Vj^��u�   �;�}�ƣ!jP�����YY�!��ujV�5!����YY�!��ujX^�3ҹ���� �R��}�!��3�^��>  �=� t�_?  �5!�����%! Yø��U��V�u��;�r"���w��+�����P������N �  Y�
�F P��`^]�U��E��}��P�����EY�H �  ]ËE�� P��`]�U��E��;�r=�w�`���+�����P����Y]Ã� P��`]�U��M�E��}�`����AP����Y]Ã� P��`]�U���V�u�M������u�E�M�L0u3�9Ut�E����   �p#E���t3�B�}� ^t�M��ap�����U��jj �uj ������]�U��} u�u�ƒ��Y]�V�u��u�u�{���Y3��MS�0��uFV�uj �5���`�؅�u^9�t@V�Q���Y��t���v�V�A���Y������    3�[^]���������`P�����Y����������`P�����Y�����U��V�u��tj�3�X��;Es�����    3��Q�u��uF3Ƀ��wVj�5��`�ȅ�u*�=� tV����Y��uЋE��t�봋E��t�    ��^]�U��V�uWV��:  Y�N�����u����� 	   �N ����  ��@t������ "   ��S3���t�^��t}�F�����N�F�����F�^�  u*������ ;�t������@;�uW�b:  Y��uV�XG  Y�F  tz�V��B��F+�H�M�F��~QRW�<  �����G�� �N�h���t���t�ϋǃ���������0�A tjSSW�{E  #����t%�N�E��3�@P�E�EPW�J<  ����;]t	�N �����E[_^]�U���  �� 3ŉE��ESV�uW�}�u������3��؍������������������������������������������������������������ɩ���p�������������������
  �@@ucP��8  Y�ȃ��t���t�у���������0�B$��
  ���t���t������������0�A$��b
  ���Z
  �3��Љ��������������������������������������
  ������������@����������	  �A�<Xw���������3�������������������������������������	  �$��3���������؉������������������������������������L	  ���� tF��t9��t/HHt���������-	  ���������	  ���������	  �����ˀ   ������*u/�������������������  ���؉�������������  ������k�
�����������������ȉ������  3��������  ��*u+������������������������r  ��������f  ������k�
�����Љ������>  ��ItE��ht8��������lt��w�,  ��   ������8lu@��   �������������� ������������ <6u�������4u�ǃ��� �  ����<3u�������2u�ǃ����������<d��  <i��  <o��  <u��  <x��  <X��  3��������3�������������P��P�*  YY��t8������P�������������  ���������A���������������b  ������P�������������  ����  ����d��  �Q  ��S��   t|��AtHHtVHHtHH�  �� ǅ����   ��������������@�   ���������������������2  ǅ����   �  ��0  ��   ��   �������   ��0  u��   �������������������t�ʋ7����������  �S  ��u�5ǅ����   �ƅ�t3�If9t����u�+����<  ��X��  HHtp���'���HH�$  ����������  t0�G�Ph   ������P������P��B  ����tǅ����   ��G�������ǅ����   ��������  �����������t3�p��t,� ��   t�+���ǅ����   �  3ɉ������}  �5V����Y�k  ��p��  ��  ��e�Y  ��g�K�����itd��nt%��o�=  ǅ����   ��y[��   �������M�����������@  ���   �������� tf���ǅ����   �z  ��@������ǅ����
   �� �  u��   ��  �����������3��  u��guVǅ����   �J;�~������=�   ~7��]  W����Y��������������t
���������
ǅ�����   ����������������G�������������P��������������������P������������VP�5�`�Ћ�����   t!������ u������PV�5$�`��YY������gu��u������PV�5 �`��YY�>-�(�����   ������F����ǅ����   j���s�����HH��������k  j'X������ǅ����   ���|���Qƅ����0������ǅ����   �^�����3��������� t��@t�G���G����@t
�G���ȋ���O�����@t;�|;�s����߁�   �������� �  u����������y3�B�����   ������;�~�Ћ��u�������u��J�����������t=�������RPWQ��  ��0����������������9~������������������N밋������E�+�F��������   t6��t�>0t-N�������0�!��u�5���I�8 t@��u�+Ɖ����������� ��  ��@t5��   t	ƅ����-���t	ƅ����+���tƅ���� ǅ����   ������+�����������+���u������P������Wj �   ��������������������Q������P������P�  ����t��u������P������Wj0�  �������� ������t}��~y��H�������Pj�E�P��������P��������=  ����u?9�����t7������������P�������E�������P�r  ����������������u��(����������#������������Q������PV�8  ����������x#��t������P������Wj ��   ����������������tP�+���3�Y������������������������������������������� _^[t
�������ap��M�3��:����������    �M�������ɋ� L��T�U��U�B@t�z t-�Jx��M������ERP�����YY���u�E��]ËE� ]�U��V�u��~W�}W�uN�u�������?�t���_^]�U��V�uW�}��G@�Et� u
�M�E�N�& S�]��~@�EP�EW� PK�K����E���E�8�u�>*uPWj?�/����E����˃> u�E�[_^]Ã%! ����������������Q�L$+ȃ����Y�;  Q�L$+ȃ����Y�;  S��QQ�����U�k�l$���   �� 3ŉE��CV�s��W��|���Ht+Ht$HtHtHtHHtHuzj��   �nj�
j�j�j_Q�FPW�K;  ����uG�K��t��t��t�e����E��F����]����E��FP�FPQW��|���P�E�P��<  ����|���h��  Q�@  �>YYt�= uV����Y��u�6�?  Y�M�_3�^�҃����]��[������������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� �����������U��SVWUj j h�u�I  ]_^[��]ËL$�A   �   t2�D$�H�3������U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�hd�5    �� 3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �yu�Q�R9Qu�   �SQ� �SQ� �L$�K�C�kUQPXY]Y[� ���U��V�u����   �F;DtP�m���Y�F;HtP�[���Y�F;LtP�I���Y�F;PtP�7���Y�F;TtP�%���Y�F ;XtP����Y�F$;\tP����Y�F8;ptP����Y�F<;ttP����Y�F@;xtP����Y�FD;|tP���Y�FH;�tP���Y�FL;�tP���Y^]�U��V�u��tY�;8tP�v��Y�F;<tP�d��Y�F;@tP�R��Y�F0;htP�@��Y�F4;ltP�.��Y^]�U��V�u���n  �v����v����v����v��~���v��~���v��~���6��~���v ��~���v$��~���v(��~���v,��~���v0�~���v4�~���v�~���v8�~���v<�~����@�v@�~���vD�~���vH�~���vL�y~���vP�q~���vT�i~���vX�a~���v\�Y~���v`�Q~���vd�I~���vh�A~���vl�9~���vp�1~���vt�)~���vx�!~���v|�~����@���   �~�����   � ~�����   ��}�����   ��}�����   ��}�����   ��}�����   ��}�����   �}�����   �}�����   �}�����   �}�����   �}�����   �}�����   �|}�����   �q}�����   �f}����@���   �X}�����   �M}�����   �B}�����   �7}�����   �,}�����   �!}�����   �}�����   �}�����   � }�����   ��|�����   ��|�����   ��|�����   ��|�����   ��|����   �|����  �|����@��  �|����  �|����  �|����  �|����  �y|����  �n|����   �c|����$  �X|����(  �M|����,  �B|����0  �7|����4  �,|����8  �!|����<  �|����@  �|����D  � |����@��H  ��{����L  ��{����P  ��{����T  ��{����X  ��{����\  �{����`  �{����^]�U��QQ�� 3ŉE�SV�uW��~!�E��I�8 t@��u������+�H;ƍp|���M$3���u�E� �@�E$��3�9E(j ��j V�u��   PQ�D`�ȉM���u3��X  ~Kj�3�X���r?�M   ��   w���c����܅�t���  �Q�+{����Y��t	���  ���M��3ۅ�t�QSV�uj�u$�D`����   �u�j j VS�u�u�c�����������   �   �Mt,�M ����   ;���   Q�uVS�u�u�(������   ��~Bj�3�X����r6�}   ;�w�������tf���  �P�lz����Y��tQ���  ���3���t@WV�u�S�u�u���������t!3�PP9E uPP��u �uWVP�u$�t`��V�����YS�����Y�Ǎe�_^[�M�3��{����U����u�M�蹓���u(�E��u$�u �u�u�u�u�uP�������$�}� t�M��ap���U��Q�� 3ŉE��MSVW3���u�E� �@�E��3�9E WW�u���u��   PQ�D`�؅�u3��   ~A�����w9�]   =   w�i������t����  �P�1y����Y��t����  �������t��PWV�y����SV�u�uj�u�D`��t�uPV�u��`��V�����Y�Ǎe�_^[�M�3���y����U����u�M�艒���u �E��u�u�u�u�uP��������}� t�M��ap���U����M�S�u�J����]�C=   w�E苀�   �X�n�����E�M���QP�   YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�E�PQ�E�P�E�jP�A�������u8E�t�E��`p�3���E�#E�}� t�M��ap�[��jh���$�����
95�
t*j����Y�e� Vh�
�S���YY��
�E������   �-����j�����Y�U����u�M��J����E��M���   �H% �  �}� t�M��ap���U��j �u����YY]�U���D�� 3ŉE��MS�A
��% �  �E��A�E��A�E�����  V���?  W�}��3ۉ}��U��E������u%���9\��u@��|��  3��}𫫫j[�  ���u��}�H��H�U܉E̋��j�^#�����]ԉUā�  �yI���A+�3�@����j����u�^�D����   �����ЅD���9\��u
B;�|��   �E̙jY#�ЋE���%  �yH���@+�3�@��j��]�_�EȋD���M�ȉM�;ȋE؋�r;E�s3�A�M�J�D��x.��t'�D���ˍx;��]ԉ}؋�r��s3�A�M�J�D��yՃ���MЋUċ���!D���B;�}�}��΍<�+�3�����M�9]�tA����+�;�}3��}𫫫������;��  +U܍u�UЋ�}�������EċEХ%  �yH���@�EЃ���ǋ}Ћ���j �]��ЉE�X+�j�E�^�T����#E؋���M���U�C�T��E�;�|ߋE����U�j+ЋE�3�Y���;�|��D���E���\����Iy�M�A���������Uԁ�  �yI���AjX+��EЋM�3�@���D����   �����ЅD���9\��uB;�|��v�}̋ǙjY#������  �yO���G�D��+�3�G��j��ˉ}���}�;��E�_r;E�s3�AJ�D��x(��t!�D���ˍx;��}���r��s3�AJ�D��yۃ���MЋUԋ���!D��B;�}�}��΍<�+�3������A���������E؁�  �yI���A�M����j �]��]�Y+��׉ẺM܋T������M�#�U��T���M����E��E�@�E�;�|׋u؋����U�j+�Y3�;�|��D����\����Iy������;���   ��3��}𫫫�M�   ����������É�  �yI���A�����j X+��M��׉]��E؋T������M�#���U��MȉT��C�E�;�|ߋű����U�j+�Y3�;�|��D����\����Iy�5�5�3�C�   �5��e���������������uȉE؁�  �yI���A��j �]���X��+ÉM��׉E܋T������M�#���U�F�T��E���|ߋ}؋uȋ����U�j+�Y3�;�|��D����\����Iy�}�jX+��ȋE������%   ��u���@u
�E�w���� u�7�M�_^��3�[��r����U���D�� 3ŉE��MS�A
��% �  �E��A�E��A�E�����  V���?  W�}��3ۉ}��U��E������u%���9\��u@��|��  3��}𫫫j[�  ���u��}�H��H�U܉E̋��j�^#�����]ԉUā�  �yI���A+�3�@����j����u�^�D����   �����ЅD���9\��u
B;�|��   �E̙jY#�ЋE���%  �yH���@+�3�@��j��]�_�EȋD���M�ȉM�;ȋE؋�r;E�s3�A�M�J�D��x.��t'�D���ˍx;��]ԉ}؋�r��s3�A�M�J�D��yՃ���MЋUċ���!D���B;�}�}��΍<�+�3�����M�9]�tA����+�;�}3��}𫫫������;��  +U܍u�UЋ�}�������EċEХ%  �yH���@�EЃ���ǋ}Ћ���j �]��ЉE�X+�j�E�^�T����#E؋���M���U�C�T��E�;�|ߋE����U�j+ЋE�3�Y���;�|��D���E���\����Iy�M�A���������Uԁ�  �yI���AjX+��EЋM�3�@���D����   �����ЅD���9\��uB;�|��v�}̋ǙjY#������  �yO���G�D��+�3�G��j��ˉ}���}�;��E�_r;E�s3�AJ�D��x(��t!�D���ˍx;��}���r��s3�AJ�D��yۃ���MЋUԋ���!D��B;�}�}��΍<�+�3������A���������E؁�  �yI���A�M����j �]��]�Y+��׉ẺM܋T������M�#�U��T���M����E��E�@�E�;�|׋u؋����U�j+�Y3�;�|��D����\����Iy������;���   ��3��}𫫫�M�   ����������É�  �yI���A�����j X+��M��׉]��E؋T������M�#���U��MȉT��C�E�;�|ߋű����U�j+�Y3�;�|��D����\����Iy�5�5�3�C�   �5��e���������������uȉE؁�  �yI���A��j �]���X��+ÉM��׉E܋T������M�#���U�F�T��E���|ߋ}؋uȋ����U�j+�Y3�;�|��D����\����Iy�}�jX+��ȋE������%   ��u���@u
�E�w���� u�7�M�_^��3�[�m����U���|�� 3ŉE��E�E��E�E�3�S3�@V�E���W�}��]��]��]��]��]���]�9E$u薧���    �W���3���  �M�щU���� t��	t
��
t��uA��A���{  �$��+�B�<wjXI���E$� ���   � :ujX����+tHHt����  3�@�j� �  X�U��jX�]��3�@�E��B�<v��E$� ���   � :uj묀�+t+��-t&��0t���C�3  ��E~��d���"  j�|���Ij�t����B�<�P����E$� ���   � :�R�����0�c����M���  3�@�E���0|*�E��u���9��s	��0@�G�F�A��0}�u��E���E$� ���   � :�I�����+�t�����-�k����E���3�@�E��E��E���u��0u�E��HA��0t��E��E���0|%�u���9��s��0@�GN�A��0}�u��E����+������-������C~��E�������d�������I�  3�@��0�E���	����j�/����A��E��B�<wj	������+t"HHt�������j����j���X�U������j����3�@�E���A��0t���1����   몍B�<v���0�9] t"�A��E���+t�HH�q����M��jX�}���j
XI��
�p����A3�@�E������9,k�
������P  
�A��0}���Q  ���9�A��0}�I�E��U��
�M�����  ��v�E�<|���E��M�OjAX�M���M�����  O8u
HAO8t��M��M�QP�E�P��&  �U�����y�ދE�u���uu�E���u+u��P  �,  �������  ����`����  y
�8�ރ�`9]��  3�f�M���  �΃�T���E��u�����  k�ȸ �  �M�f9r��}����M���M��M��y
�U΋�3�% �  �E���  #�#��]�����  �]ԉ]؉]܉u�f;��+  f;��"  ���  f;��  ��?  f;�w�]��  f��u$F�E�����u�u�}� u�}� u3�f�E���  f��uF�A����u�u	9Yu9t�j��_�E��U؉}��}���~\�uč4F�A�E���� �E���}����}�z��]�;z�r;}�s3�@��E��z���tf��E�����I�E�����M��}��E���@O�E��}�����u��U܋}ԁ��  �U�f��~;��x2�E؋ȋ����U��E���Ҹ��  ����}ԉU��U�f���f��i���  �f��y]�]��������E���E�tC�M؋����M��m�	E��E���������M��U܉E؉}�u�j �ۉU�[tf��3�Gf�f�Eԋ}��f�EԺ �  f;�w���� �� � u@�Eփ��u4�Eډ]փ��u f�E޹��  �]�f;�uf�U�F�f@f�E��@�EڋM��@�E֋M���  f;�sf�E�u�f�EċE؉EƉM�f�u��3�f9E���H%   � ���Ẻ]ĉ]ȋE��u����1����E��MċUƋu����23��ˋË�Ӎ_�#��  �   �j��ˋË����Ë�j�ˋ�[�}�E�f�f�G
�W�w�ËM�_^3�[�>f���Ð%k%�%�%W&�&�&V'8'�'�'b'U���   �� 3ŉE��US�]V� �  #��u3ɸ�  A#�W�]��E������E������E����?�U��E�f��t�C-��C �}f��u:����   9}��   3�f�� �  f;�����$ �C�Kf�C0 ����  f;���   �E�   �f��M;�u��t�   @uh���Gf�}� t=   �u��u0h���;�u%��u!h ��CjP�d���������  �C�h��CjP�C���������  �C3��9  �֋�i�M  ����������Hk�M����ȋE�E�3��M���f�E��ٸ���`3�f�u�}�M��E�   �E���  �E��?  ���!  y�ٸ8��`�M����
  �u��U�u��}���T�E�����  k�ȸ �  ��x���f9r��}ĥ��Mĥ�MƉ�x����y
�E�}�1E�%�  ���  �E�Ǿ �  !u��}����E�N�]��]��]�]��}�f;��J  f9u��u��=  f;}��3  f;}�w�]��<  f��u G�E�����}�u��u��u3�f�E��$  f�}� uG�A����}�u	9Yu9t�j��^�E��U�u��u���~o�u��F�q�M��E���|����8����B��]��48;��u���r;�s3�F��u��B���tf��E���|�������I�E���|��������x����u��E���@N�E��u����w����}��E��u����  �E�f��~;��x2�E�������E�E��������  ���u��E��E�f���f��q���  �f��ye�]��������3҉}��}��E�B�U�tG�M�����M��m�	E��E���������M��]��E�u�u�j �]����}�[tf��f�f�E��u��f�E� �  f;�w���� �� � u@�E���u4�E��]���u f�E����  �]�f;�uf�M�G�f@f�E��@�E��M��@�E�M���  f;�s f�E�}�f�E��E�E�u��M�U�f�}��!3�f9E���H%   � ���E��Ӊu��U�u��E��M���������U�u��E�����?  f;���  �E��ȋEڋ�3��� �  �}���  #�#ωE������  �]��]��]�]��}�f;��@  �E�f;E��3  f;}��)  f;}�w�]��2  f��u G�E�����}�u��u��u3�f�E��  f��uG�E�����}�u�}� u�}� t���j�U��M�X����~X�}��E؍<W�E��}����ЋA��]��<;�r;�s3�@��E��y���tf��}��E�����N�}��E�����U��E���BH�U��E�����}��u����  f����   �]��]���x,�E�ȋ����E�������  ����]��u�f��Љ]��U�j [f��~[f�M� �  f;�w���� �� � ��   �E�����   �E��]�����   f�E����  �]�f;�u|� �  f�E�G�|�U���  �f��y���������}��}��E��E�tG�]�ˋ��������������M��]�U�u�j ���}��u�[�M���3�f��@f�f�M��U��<���f@f�E��@�E��u��@�E��  f;�s f�E�}�f�E��E�E�u�U�u�f�}��3�f9E���H%   � ���E����E�M��E��}f�t6���}���/3�f�� �  f9E�����$ �A3�@�A�A0�Y�  �}�jX;�~�E��}������?  3�j�}�f�E�]�_�ʋ���������Љu��]�Ou�}�j �]��U�u�[��y7�߁��   ~-�]��ʋ�������������O�]�u����]��U�u�3ۋu��E��~@�ω}��M��E�����   �u��}ĥ���}��ʋ����ЋE����4 ���ǋ������ЋE����8�M�;�r;�s�B��;�r��s3�A�ɋM���tF�Eȍ<;�r;�sF�U�u�ҋ����U��U��?Ћ����6��M��E���0��E�AH�U�M��]�E���~�E�E��>����u��}��A���<5|C�	�99u�0I;�s�;�sAf���E�*Ȁ��H�Ɉ\3�@�M�_^3�[�\���À90uI;�s�;�s΋M�3�f�� �  f9E�����$ �A3�@�A�0����3�SSSSS�}����U��M3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tƋѻ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t;�u �  ]Ã�@]�@�  ]�U�����}�f�E�3ɨtjY�t���t���t��� t���t��   SV���ֻ   W�   #�t&��   t��   t;�u��   �
����   ��   t;�u��   ���   ���   ��t��   �}�E����#�#��;���   V�=  ��Y�E��m���}��E�3��tj^�t���t���t��� t���t��   �Ћ�#�t*��   t��   t;�u��   ���   ���   ��   t��   u��   ���   �   ��t��   �=���  ���]�E�3Ʉ�yjY�   t���   t���   t����t���   t��   �л `  #�t*��    t�� @  t;�u��   ���   ���   j@%@�  [+�t-�  t+�u��   ���   ���   ��#}��#��;���   P�$���P�E�\  YY�]�E3Ʉ�yjY�   t���   t���   t���   t���   t��   �п `  #�t*��    t�� @  t;�u��   ���   ���   %@�  +�t-�  t+�u��   ���   ���   ��3�Ω t��   ������_^[��U��M3���t@��t����t����t����t�� ��   t��V�Ѿ   W�   #�t#��   t;�t;�u   �   �   �с�   t��   u���_^��   t   ]�U��E��u�Q����    �������]Ë@]�U��M���u�,���� 	   �8��x$;�1s������������D��@]������� 	   踘��3�]�U��V�u��u	V�   Y�/V�,   Y��t�����F @  tV�U���P�D  Y��Y��3�^]�U��SV�u3ۋF$<uB�F  t9W�>+~��~.W�vV����YP�  ��;�u�F��y����F��N ���_�N�f �^��[]�j�   Y�jh��� ���3��}�!}�j�n���Y!}�3��]�u�;5!��   �!����t]�@�tWPV����YY�E�   �!���@�t0��uP�����Y���tG�}����u�@tP�����Y���u	E܃e� �   F녋]�}�u�!�4�V����YY��E������   ����t�E��}���Ë]�}�j����Y�jh������3��}�j荩��Y!}�j^�u�;5!}S�!����tD�@�tP��  Y���tG�}��|)�!���� P�T`�!�4��,T��Y�!�$� F��E������   ���ݍ��Ë}�j�n���Y�jh������u���u�g����  蓏��� 	   �   ����   ;5�1��   ��������������D8��tcV�  Y�e� ����D8t�u�uV�_   ������%���� 	   �����  ����}��E������
   ���)�u�}�V��  Y�躎���  ����� 	   觕����������U���  �,  �� 3ŉE��E�M3�W����@�����D�����<�����,���9Uu3���  ��u�O���!8�|����    �=�������  SV������������0������������\$�����t��u+�E�Шu����!8� ����    �����L  ��@����D tjRRP�M  ����@�������Y���  ��0�������D��   �Yz���@l3�9��   �����P��0���������4��@�����`����  9�@���t����  ��`��D���!�$����ʉ������4���9}�~  3���8���ǅ���
   ����  �	3���
����@�����0�������|8 t�D4�E�j�E�M��d8 P�Z��P�$���Y��tD��D�����4���+�E����  jR��<���P�  �������  ��4���@��8����&j��4�����<���P�  �������  ��4���3�QQ@��8���j��4����E�Pj��<���PQ������t`��������k  j ��$���QP�E�P��0�������4� `����  ��8���������,���9�$����!  ��@��� ��   j ��$���Pj�E�P��0����E�����4� `����  ��$�����   ��,���G�   ��t��u3�3�f;������<�����8���������4�����8�����@�����t��uU��<����`  Yf;�<����  ����@��� t$jXP��<����7  Yf;�<�����  G��,�����8�����4���;E������#��0�������G�D4����D8   ��@����  ��@����  ��0�������D��U  ��D���3���8�������   ��<���9u��  3�+�<�����H�����@���;EsD�
B@��#�����
��@�����<���u��,����CA��#������<���CA��@������  r��������H���+�j ��(���PS��H���P��0�������4� `����  �(�����D���9�(�����  ��<���+�;E��<����5����  �ʀ���   ��@���9u��  ǅ���
   ����� ��,�����+������H���;Es>�1������@���f;����ujYf���@���������f�3�������  r��������H���+�j ��(���PS��H���P��0�����,�������4� `��8�����<�������  �(�����D�����<���9�(�����  ��@�����+�;E� ����  �]��$�������  ǅ���
   ����� ��$���+ʋ������H���;�s;�>������$���f;����uj^f�0��$�������f�8�������  r�3�VVhU  ������Q��H���+��+���P��PVh��  �t`��8�����<�����4�������   3ɉ�@���j +���(���RP������������P��0�������4� `��t��@����(�����4�����@���;����`��@�������4�����8���;�Q��$�����D�����+���<���;�������7j ��(���Q�u��D����4� `��t
��(���3���`����D�����uc��t$j[;�u����� 	   �ӆ����?V�܆��Y�6��0������������D@t	�:u3�� �҆���    蓆���  ����+�,�����^[�M�3�_�QL����jh(��s�������u؉u܋}���u�R����  �~���� 	   �   ����   ;=�1��   �����E�߃�������D��tpW�  Y�e� �E����Dt�u�u�uW�g   ������������ 	   �ƅ���  �މu؉]��E������   ���+�}�]܋u�W�  Y�蕅���  ������ 	   肌���֋��Ƀ���U��QQV�uWV�  ���Y;�u菅��� 	   �ǋ��D�u�M�Q�u�uP��`��u�`P�>���Y�Ӌ�����������d0��E��U�_^��U���� V�   V�&���Y�M�A��t	�I�q��I�A�A�A   �A�a �^]Ë� ��3�9!���U���S�]W�}��u��t�E��t�  3���E��t��V�����v褄��j^�0�f����X�u�M���b���E�3�9��   u`f�E��   f;�v9��t��tWVS�yI�����Z���� *   �O����0�}� t�M��ap���^_[�Å�t��t_��E��t��    �ӍMQVWSj�MQV�u�p�t`�ȅ�t9uu��E��t����`��zu���t��tWVS��H�����̓��j"^�0菊���q���U��j �u�u�u�u�������]�����������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ��U���S�]V�����t�Etj�  Y����  ��t�Etj�  Y����u  ����   �E��   j�]  �EY�   #�tT=   t7=   t;�ub��M�������{L�H��M�����{,���2��M�����z�����M�����z�������������   ����   �E��   W3���tG�M���������D��   ��EPQQ�$�  �E�U��� ������E=����}3���G�W��3�����AuB�E�����f�E��E����;�})+ȋE��E�t��uG���E��E�t   ��E��m�Iu��E��t���E��3�G��_tj�  Y�����t�E tj ��  Y���3���^��[��U��j �u�u�u�u�u�u�   ��]�U��E3ɉH�ES�H�E3ۉH�MCW��t�E��  �	X��}��t�E��  ��H��t�E��  ��H��t�E��  ��H��t�E��  ��H�MV�u�����3A��1A��M���3A��1A��M����3A��1A��M����3A��1A��M����3A#�1A�9  ����t�M�I��t�E�H��t�E�H��t�E�H�� t�E	X��   #�t5=   t"=   t;�u)�E��!�M���������M��������E� ���   #�t =   t;�u"�E� ���M�������M�������E�M��3���� 1�E	X �}  t,�E�` �E� �E�X�E	X`�E�]�``�E��XP�:�M�A �����A �E� �E�X�E	X`�M�]�A`�����A`��E�XP�f  �EPjj W��`�M�At�&��At�&��At�&��At�&��At�&ߋ��������� t/HtHtHu(�   � �%����   ���%����   ��!������� tHtHu!��#�   �	�#�   ��}  ^t�AP���AP�_[]�U��E��t�����w�t~��� "   ]��g~��� !   ]�jhH��*|���=�|[�E�@tJ�=� tA�e� �U�.�E� �8  �t�8  �t3��3�@Ëe�%� �e��U�E������
�࿉E�U�|���U��Q�}����E���U��Q��}��M�E#E��f#M�f����E�m�E���U��QQ�M��t
�-��]���t����-��]�������t
�-��]����t	�������؛�� t���]����U��Q��}��E���U���S�]3�V�N@  W�E���S�S9U�@  �ʉM�U��U�U��}䥥��u��}������������ҋ��������E�������3ɉ�s�{�E;�r;E�s3�A���t��3ɍp;�r��s3�A�s��tG�{�U�3���M�;�r;�s3�@�K��tG�{�U}�u�e� ���������?��M҉�s�C�9�u��:�E�}�M;�r;�s3�B��U����t'�N3�;�r��s3�B��K�M�u���t@�E�C�C�EH�E�s�E��������N@  3�9Su.�S��������ЋE�������  ��E���tۉS�s�S�� �  u4�;�s���������E�������  ��E��� �  tى;�s�S_^f�C
[��jhh��6y���}���u�R{��� 	   �   ����   ;=�1��   �����E��߃�������D��ttW�j  Y3��u��E�����Dt(W�_  YP��`��u�`���u��t�z���0��z��� 	   ����u��E������
   ���!�}�u�W�w  Y��z��� 	   �Z�������x���U��V�uW�����u�qz���    �2�����E�F�t9V����V���-  V�����P�  ����y�����~ t�v�s>���f Y�f ��_^]�jh����w������}�3��u������u��y���    赀������w����F@t�f ��V�9���Y�e� V�?���Y���}��E������   �ǋu�}�V�}���Y�jh���mw���}����������4���~ u0j
�ƒ��Y�e� �~ uh�  �FP�P`�F�E������*   ��������������P��`3�@�?w��Ë}j
�Г��Y�U��EVW��x`;�1sX��������������Dt=�<�t7�=Pu3�+�tHtHuQj��Qj��Qj���`�����3���x��� 	   �fx���  ���_^]�U��M���u�Lx���  �xx��� 	   �B��x&;�1s������������Dt�]��x���  �9x��� 	   ��~�����]�U��M��������������P��`]�U���SV�u��t�]��t�> u�E��t3�f�3�^[��W�u�M��V���E����    u�M��t�f�3�G�   �E�P�P����YY��t@�}��t~';_t|%3�9E��P�u�wtVj	�w�D`�}���u;_tr.�~ t(�t�13�9E��3�GP�u�E�WVj	�p�D`��u�.w������ *   �}� t�M��ap���_�6���U��j �u�u�u�������]�U��Q�����u
�  �����u���  ��j �M�Qj�MQP��`��t�f�E��U���EW��������Dz	��3��   Vf�u�Ʃ�  u|�M�U���� u��tj�ٿ�������Au3�@�3��EuɉM��y���M�O�Et�f�u�U���  f#�f�u��t� �  f�f�u�Ej QQ�$�1   ���#j ��QQ�$�   �������  �����  ^�E�8_]�U��QQ�M�E�E�]����  ��%�  �f�M��E���̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� jh���Ps���u���u�8u���  �du��� 	   �   ��xy;5�1sq��������������D8��tSV����Y�e� ����D8tV�U   Y����u��� 	   ����}��E������
   ���)�u�}�V����Y��t���  ��t��� 	   �{�������r���U��VW�}W����Y���tP����u	���   u��u�@Dtj�����j�������YY;�tW�����YP��`��u
�`���3�W�9���Y������������D9 ��tV�t��Y����3�_^]�U��V�u�F�t �Ft�v�Q8���f����3�Y��F�F^]á����t���tP��`�3�PPjPjh   @h����`����%(`�%�`������h�X�@��Y����̃=  uK����t�Q�@<�@�Ѓ���    V�5��t���p���V������    ^�                                                                                                                                                                                                                           �  � 0� B� X� h� t� �� �� �� �� �� �� �� � � 2� D� Z� l� z� �� �� �� �� �� � ,� F� `� v� �� �� �� �� �� ��  � 
� � &� :� F� \� n� ~� �� �� �� �� �� �� �� �� � � .� @� T� f� z� �� �� ��         �X        d���)���3�        xX��                        `�
R       �   H� H�     `�
R          �� �� ���Q��?      @�������?�������?�������?ffffff�?��Q��?�������N���������������C-DT�!	@-DT�!�?�� a  � p� � � �� ` �a � � � ` � P� `� p� �� � �� �% �� & �a tool_AMa_1D_Snap        d:\applications\maxon\cinema 4d r14 demo\plugins\ama_1d_snap\source\ama_1d_snap.cpp     AMa_1D_Snap.tif ���Q��?�������?�������?��Q��?�������?ffffff�?      �?      @      B@���������������������N���������������C-DT�!	@-DT�!�?COMMANDLINE number of arguments:    --help  -help   -SDK is here :-)   -SDK    -SDK executed:-)   -plugincrash    C4DSDK - Edit Image Hook:   ��pn �������N���������������C-DT�!	@-DT�!�?res     �������N���������������C-DT�!	@-DT�!�?d:\applications\maxon\cinema 4d r14 demo\resource\_api\c4d_general.h       %s  �������N���������������C-DT�!	@-DT�!�?���� @�     d:\applications\maxon\cinema 4d r14 demo\resource\_api\c4d_baseobject.cpp       ����MbP?d:\applications\maxon\cinema 4d r14 demo\resource\_api\c4d_resource.cpp #   M_EDITOR    �������N���������������C-DT�!	@-DT�!�?�������N���������������C-DT�!	@-DT�!�?�������N���������������C-DT�!	@-DT�!�?d:\applications\maxon\cinema 4d r14 demo\resource\_api\c4d_file.cpp     �������N���������������C-DT�!	@-DT�!�?d:\applications\maxon\cinema 4d r14 demo\resource\_api\c4d_basebitmap.cpp       d:\applications\maxon\cinema 4d r14 demo\resource\_api\c4d_misc\datastructures\basearray.h      d:\applications\maxon\cinema 4d r14 demo\resource\_api\c4d_libs\lib_ngon.cpp          �?�������������d:\applications\maxon\cinema 4d r14 demo\resource\_api\c4d_pmain.cpp                  �      ���������������-DT�!�?-DT�!��RUUUUU�?        v�F�$I�?������ɿ��3Y�E�?#Y��q���n����?��;
9��� ��/I�?hK����d��?81�U����H!G�?��#�$�����0|f?�K�RVn���TUUUU�?        ~I�$I�?g����ɿHB�;E�?����q���{雮?�x��֚��                   �      �?       @       @      �?      �?      @>��1|�MC                                            �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������                                      �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      �D�V�u�    R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
       R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
   R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
     R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
   R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
         R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
       R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
         R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
         R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
     R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
         R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
     R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
     R 6 0 3 4  
 -   i n c o n s i s t e n t   o n e x i t   b e g i n - e n d   v a r i a b l e s  
     D O M A I N   e r r o r  
     S I N G   e r r o r  
     T L O S S   e r r o r  
    
     r u n t i m e   e r r o r          ��   pz	   �z
    {   h{   �{    |   h|   �|   0}   �}   �}   `~   �~   �~    �!    �"   �x   x�y   ��z   ���   Ђ�   ؂R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
     R u n t i m e   E r r o r ! 
 
 P r o g r a m :     < p r o g r a m   n a m e   u n k n o w n >     . . .   
 
     M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y               �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��log log10   exp pow asin    acos    exp10   atan    ceil    floor   modf    sin cos tan sqrt       �U��?�wB%�K�=      �?   �[��?(�6N�g�=      �?   $�?V�`t� >      �?   ��տ?��2n{a>      �?   ����?��M��=      �?   H{��?{4�r>      �?   Pא�?"�"�>      �?   �u[�?��*��>      �?   ����?G�0��_(>      �?   4wb�?��i^^?(>      �?   ��0�?p3���>      �?   @��?F��M>      �?   8M��?�B�V��>      �?   ��d�?}B��a.>      �?   ȴ�?d�����>      �?   g��?�ߊ��>      �?   �@�?�f\���*>      �?   �~e�?�-��f>      �?   �]%�?D	�G��?>      �?   ���?�\����>>      �?   X���?�1��#>      �?   �E�?��h��>      �?   �?��?�ⳇ��>      �?   ����?�$	�49>      �?   x�8�?k���0H<>      �?   ����?r��ش8>      �?   8fm�?�"m>">      �?   ħ �?[��<c�'>      �?   �k��?"���%>      �?   ���?݉@fR�8>      �?   ����?��T���:>      �?   T�!�?3&�F>      �?   � ��?<����[#>     ��?   �%�?�Y:/(A6>      �?   ����?��N��2>     ��?   8O�?�r�!'	>      �?   ��r�?���8{K>     ��?   �p��?9��l�9$>      �?   �
G�?�aj	�i9>     ��?   T|��?'\�|#<>      �?   $��?�}�dj�#>     ��?   �Wn�?׈MVx:>      �?   ,���?1�8o,>     ��?   D�$�?	c�/�
>      �?   @ |�?��x7|�1>     ��?   |���?��9>      �?   p #�?�IA��u=>     ��?   �s�?�x ٴ4>      �?   p���?edf�&�.>     ��?   ,�?��f���A>      �?   h�*�?v����2>     ��?   $gN�?RE\��K>      �?   �q�?'^��IE>     ��?   DΒ�?��&a��H>      �?   L���?�&KrQF>     ��?   ,���?�#/�'�>      �?   إ��?]X�c�?>     ��?    ��?�Ԯ}�>      �?   �e.�?�IdW�A>     ��?   �K�?���ΐ?>      �?   Xg�?��4*�A>     ��?   _��?�[�ǆJ>      �?   ���?1���0H>     ��?   ���?�hc#�]G>       @   ,*��?�Q�x
�F>     @ @   p���?ek�R�.N>     � @   �� �?�Ӿ�n@>     � @   �b�?�����O>      @   $Q/�?CJ���O>     @@   ��E�?������G>     �@   �[�?�3E�{A>     �@   T�p�?�SfI�S:>      @   X΅�?B6)�1�<>     @@   �3��?>ځ���7>     �@   $��?s(��N>     �@   @���?V�
6�f=>      @   (���?��{��>     @@   (W��?��-�Jg >     �@   ����?��"a�PK>     �@   xm�?,S��ڤ6>      @   ���?�6��hb">     @@    �-�?�k,�<>     �@   X�>�?�0����=>     �@   �O�?�׀IX�H>      @   �-_�?���
@>     @@   ��n�?���2E>     �@   �P~�?�=�ő�8>     �@   lj��?�[j&,>      @   L7��?��x��82>     @@   ����?c�#V�B>     �@   0��?7ڨ.�Y>     �@   P���?�[�p&>      @   ؔ��?h4�M��A>     @@   � ��?E�p�l E>     �@   �+��?�o�$�E>     �@   h��?\���*�K>      @   ���?-�?��B>     @@   P8�?�(l�|�@>     �@   �p!�?u���@�J>     �@   @p-�?�V��1>      	@   �89�?����5>     @	@   <�D�?��ƀ�7>     �	@   h)P�?R`D�OG>     �	@   �T[�?9%� ��K>      
@   �Mf�?��/�<>     @
@   �q�?�Ò��?>     �
@   �{�?4��2G<>     �
@   L��?Â���|/>      @   �Y��?���s�
@>     @@   �k��?��Ò�a@>     �@   XS��?x(3��u8>     �@   ���?v�O,ib>      @   ȥ��?�&L͒C>     @@   ���?��}��L>     �@   �X��?Lo����>     �@   �x��?-�Ϡ�9>      @   �s��?6FID?9>     @@   8J��?����gsL>     �@   d���?��y>     �@   ���?>�&�09C>      @   ����?
��<�A>     @@   (J�?I�V	C>     �@   `w�?��^@�N>     �@   ���?�#��%�@>      @   �s�? �M�K>     @@    D'�?ή�Q��->     �@   ��.�?9!���G>     �@   ��6�?.����1>      @   >�?.1�NcB>      @   �cE�?�sǔ�1>     @@   L�L�?�n�HN>     `@   H�S�?�W��$>     �@   8�Z�?
Ȃ�q�;>     �@   ��a�?N�/�[7>     �@   (�h�?�=�mC>     �@   0oo�?�H75M>      @   Hv�?P��.�#>      @   �|�?�G���7>     @@   �*��?�#4��2I>     `@   ����?o���oJ>     �@   ����?���-��#>     �@   ���?�h��%F>     �@   @��?R�x^D>     �@   PP��?�� s�@>      @   4L��?P�_!
�#>      @   4��?��:#�G>     @@   L��?qg�:&J>     `@   Hɹ�?5L$.��4>     �@   \w��?!�1�C>     �@   ���?���[<>     �@   D���?��<���=     �@   ���?��
~���=      @   �y��?������B>      @   ����?�~.���4>     @@   h��?��u�|�8>     `@   �E��?A8yL;>     �@   �h��?��41��C>     �@   �{��?-���+oF>     �@   $��?x���O>     �@   s��?�՝m�T2>      @   �W��?����=>      @   �-�?î�\�=>     @@   ��?���\=�=     `@   ��?j\&">     �@   �X�?��1�D>>     �@   ���?�#O#`�I>     �@   ��?�}���0>     �@   ��?���F\IE>      @   t{#�?��ׯ,B>      @   0�'�?�E� ]�$>     @@   ,>,�?��ކ?5>     `@   ��0�?��iIqE>     �@   ��4�?�ha�;>     �@   �9�?��A���D>     �@   �.=�?̤KF�w�=     �@   DMA�?�����=      @   `E�?ap�I0�H>      @   �gI�?��:���->     @@   �cM�?��%Q>     `@   @UQ�?Ly5ښoE>     �@   �;U�?v�g�0�/>     �@   �Y�?jv�U�G>     �@   �\�?�����yK>     �@   ,�`�?A%My��>      @   md�?���H>      @    h�?�p���M>     @@   0�k�?k��}<>     `@   �ho�?����f7O>     �@   ��r�?���}�O>     �@    �v�?+��i�I>     �@   @z�?�b�B'=>>     �@   `�}�?Z����M>      @   ����?1�����M>      @   �a��?R�~���=     @@   t���?QNT	��B>     `@   x��?�W3c�L>     �@   g��?�+(����=     �@   D���?q���J�K>     �@   L��?� ;,*>     �@   8!��?������D>      @   ,O��?� ����E>      @   Du��?��in]D>     @@   ����?%����3F>     `@   P���?^��F"VM>     �@   ����?�}�30}->     �@   @���?�~F	y�;>     �@   ����?l	R(>     �@   躰�?��\�7`>      @    ���?�dg���;>      @   ���?�;Sv�@E>     @@   <|��?�����M>     `@   �Y��?|}�;�2>     �@   ,0��?�<v��G>     �@   $ ��?̯�/p�">     �@   ����?���\(0>     �@   |���?[s$���F>      @   I��?�d�ӔV>      @   T���?���0)LK>     @@   h���?�)�5G�5>     `@   XY��?�|��zJ>     �@   @���?W�޾�L?>     �@   0���?����6:>     �@   <3��?��Q���B>     �@   x���?7o��/�M>      @   �Q��?�Kc�Z�0>      @   ����?�z-�A5>     @@   Z��?"B�DcI>     `@   ����?��`I�.>     �@    L��?L�d�%>     �@   ���?"�l"w �=     �@   �(��?�?��!>     �@   ���?��j^�J>      @   8���? ϞH��0>      @   LL��?���%�C>     @@   T���?��J�+N>     `@   d���?;l�>�0>     �@   �B��?�^{v�@>     �@   Ȋ��?�@Y˕B>     �@   @� �?T�l���0>     �@   ��?w4n4>      @    G�?�oN�=�;>      @   h|�?�L�{�/>     @@   <�	�?B�nu5>     `@   ���?���`�,+>     �@   d�?����5>     �@   �$�?l��  >     �@   �C�?~+^��M>     �@   �^�?�PK�QD >      @   ,u�?^{�#tF>      @   |��?�^4K�� >     @@   ���?��4�O
>>     `@   ���?XEړ� J>     �@   ���?(�gԹ�,>     �@   �� �?43-spF>     �@   ��"�?P`E5�+*>     �@   ��$�?=�QQ�D>       @-DT�!�?\3&��<e+000     �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          �      	   m s c o r e e . d l l   CorExitProcess  k e r n e l 3 2 . d l l     FlsAlloc    FlsFree FlsGetValue FlsSetValue InitializeCriticalSectionEx CreateSemaphoreExW  SetThreadStackGuarantee CreateThreadpoolTimer   SetThreadpoolTimer  WaitForThreadpoolTimerCallbacks CloseThreadpoolTimer    CreateThreadpoolWait    SetThreadpoolWait   CloseThreadpoolWait FlushProcessWriteBuffers    FreeLibraryWhenCallbackReturns  GetCurrentProcessorNumber   GetLogicalProcessorInformation  CreateSymbolicLinkW SetDefaultDllDirectories    EnumSystemLocalesEx CompareStringEx GetDateFormatEx GetLocaleInfoEx GetTimeFormatEx GetUserDefaultLocaleName    IsValidLocaleName   LCMapStringEx   GetCurrentPackageId �8U S E R 3 2 . D L L     MessageBoxW GetActiveWindow GetLastActivePopup  GetUserObjectInformationW   GetProcessWindowStation    ��   ȯ   Я   د   �   �   ��    �	   �
   �   �    �   (�   0�   8�   @�   H�   P�   X�   `�   h�   p�   x�   ��   ��   ��   ��   ��   ��   ��    ��!   ��"   Ȱ#   а$   ذ%   �&   �'   �)   ��*    �+   �,   �-   �/    �6   (�7   0�8   8�9   @�>   H�?   P�@   X�A   `�C   h�D   p�F   x�G   ��I   ��J   ��K   ��N   ��O   ��P   ��V   ��W   ��Z   ȱe   б   ر  ܱ  �  ��   �  �  �  $�  0�	  <�  H�  T�  `�  l�  x�  ��  ��  ��  ��  ��  ��  ̲  ز  �  �  ��  �  �   �  ,�   8�!  D�"  P�#  \�$  h�%  t�&  ��'  ��)  ��*  ��+  ��,  ��-  Գ/  �2  �4  ��5  �6  �7  �8  (�9  4�:  @�;  L�>  X�?  d�@  p�A  |�C  ��D  ��E  ��F  ��G  ĴI  дJ  ܴK  �L  ��N   �O  �P  �R  $�V  0�W  <�Z  L�e  \�k  l�l  |��  ��  ��  ��  ��	  ��
  ĵ  е  ܵ  �  ��   �  �  $�,  0�;  H�>  T�C  `�k  x�  ��  ��  ��	  ��
  ��  Ķ  ж;  �k  ��  �  �  �	  (�
  4�  @�  L�;  X�  h�  t�  ��	  ��
  ��  ��  ��;  ȷ  ط	  �
  �  ��  �;   �  0�	  <�
  H�  T�;  l�   |�	   ��
   ��;   ��$  ��	$  ��
$  ȸ;$  Ը(  �	(  �
(  ��,  �	,  �
,   �0  ,�	0  8�
0  D�4  P�	4  \�
4  h�8  t�
8  ��<  ��
<  ��@  ��
@  ��
D  ��
H  ȹ
L  Թ
P  �|  �|  ��رB   (�,   �q   ��    ��   ��   (��   4��   @��   L��   X��   d��   p��   |��   ���   ���   ��C   ���   ���   ĺ�   �)   к�   �k   а!    �c   ȯ   �D   �}   $��   Я   <�E   �   H�G   T��   �   `�H   ��   l��   x��   ��I   ���   ���   бA   ���    �   ��J   �   Ļ�   л�   ܻ�   ��   ���    ��   ��   ��   $��   0��   <�K   H��   T��   �	   `��   l��   x��   ���   ���   ���   ���   ���   ���   ̼�   ؼ�   ��   ��   ���   ��   ��    ��   ,��   8��   �#   D�e   �*   P�l   ��&   \�h   �
   h�L   8�.   t�s    �   ���   ���   ���   ��M   ���   ���   ��>   Ƚ�   ��7   Խ   (�   �N   @�/   �t   ��   ���   �Z   0�   �O   �(   �j   ��   (�a   8�   4�P   @�   @��   L�Q   H�   X�R   0�-   d�r   P�1   p�x   ��:   |��   P�   ��?   ���   ��S   X�2   ��y   �%   ��g   �$   ��f   Ⱦ�    �+   Ծm   ��   ��=   ��   ��;   ���   H�0   ��   �w   �u   (�U   X�   4��   @�T   L��   `�   X��   x�6   d�~   h�   p�V   p�   |�W   ���   ���   ���   ���   x�   ĿX   ��   пY   ��<   ܿ�   ��   ��v    ��   ��   �[   ذ"   �d   $��   4��   D��   T��   d��   t��   ��   ��\   ���   ���   ���   ���   ���   ��   ���   ��]   `�3   �z   ȱ@   ��   ��8   $��   ��9   0��   ��   <�^   H�n   ��   T�_   p�5   `�|   Ȱ    l�b   ��   x�`   h�4   ���   ��{    �'   ��i   ��o   ��   ���   ���   ���   ��   ��   �F   (�p   a r     b g     c a     z h - C H S     c s     d a     d e     e l     e n     e s     f i     f r     h e     h u     i s     i t     j a     k o     n l     n o     p l     p t     r o     r u     h r     s k     s q     s v     t h     t r     u r     i d     u k     b e     s l     e t     l v     l t     f a     v i     h y     a z     e u     m k     a f     k a     f o     h i     m s     k k     k y     s w     u z     t t     p a     g u     t a     t e     k n     m r     s a     m n     g l     k o k   s y r   d i v       a r - S A   b g - B G   c a - E S   z h - T W   c s - C Z   d a - D K   d e - D E   e l - G R   e n - U S   f i - F I   f r - F R   h e - I L   h u - H U   i s - I S   i t - I T   j a - J P   k o - K R   n l - N L   n b - N O   p l - P L   p t - B R   r o - R O   r u - R U   h r - H R   s k - S K   s q - A L   s v - S E   t h - T H   t r - T R   u r - P K   i d - I D   u k - U A   b e - B Y   s l - S I   e t - E E   l v - L V   l t - L T   f a - I R   v i - V N   h y - A M   a z - A Z - L a t n     e u - E S   m k - M K   t n - Z A   x h - Z A   z u - Z A   a f - Z A   k a - G E   f o - F O   h i - I N   m t - M T   s e - N O   m s - M Y   k k - K Z   k y - K G   s w - K E   u z - U Z - L a t n     t t - R U   b n - I N   p a - I N   g u - I N   t a - I N   t e - I N   k n - I N   m l - I N   m r - I N   s a - I N   m n - M N   c y - G B   g l - E S   k o k - I N     s y r - S Y     d i v - M V     q u z - B O     n s - Z A   m i - N Z   a r - I Q   z h - C N   d e - C H   e n - G B   e s - M X   f r - B E   i t - C H   n l - B E   n n - N O   p t - P T   s r - S P - L a t n     s v - F I   a z - A Z - C y r l     s e - S E   m s - B N   u z - U Z - C y r l     q u z - E C     a r - E G   z h - H K   d e - A T   e n - A U   e s - E S   f r - C A   s r - S P - C y r l     s e - F I   q u z - P E     a r - L Y   z h - S G   d e - L U   e n - C A   e s - G T   f r - C H   h r - B A   s m j - N O     a r - D Z   z h - M O   d e - L I   e n - N Z   e s - C R   f r - L U   b s - B A - L a t n     s m j - S E     a r - M A   e n - I E   e s - P A   f r - M C   s r - B A - L a t n     s m a - N O     a r - T N   e n - Z A   e s - D O   s r - B A - C y r l     s m a - S E     a r - O M   e n - J M   e s - V E   s m s - F I     a r - Y E   e n - C B   e s - C O   s m n - F I     a r - S Y   e n - B Z   e s - P E   a r - J O   e n - T T   e s - A R   a r - L B   e n - Z W   e s - E C   a r - K W   e n - P H   e s - C L   a r - A E   e s - U Y   a r - B H   e s - P Y   a r - Q A   e s - B O   e s - S V   e s - H N   e s - N I   e s - P R   z h - C H T     s r     a f - z a   a r - a e   a r - b h   a r - d z   a r - e g   a r - i q   a r - j o   a r - k w   a r - l b   a r - l y   a r - m a   a r - o m   a r - q a   a r - s a   a r - s y   a r - t n   a r - y e   a z - a z - c y r l     a z - a z - l a t n     b e - b y   b g - b g   b n - i n   b s - b a - l a t n     c a - e s   c s - c z   c y - g b   d a - d k   d e - a t   d e - c h   d e - d e   d e - l i   d e - l u   d i v - m v     e l - g r   e n - a u   e n - b z   e n - c a   e n - c b   e n - g b   e n - i e   e n - j m   e n - n z   e n - p h   e n - t t   e n - u s   e n - z a   e n - z w   e s - a r   e s - b o   e s - c l   e s - c o   e s - c r   e s - d o   e s - e c   e s - e s   e s - g t   e s - h n   e s - m x   e s - n i   e s - p a   e s - p e   e s - p r   e s - p y   e s - s v   e s - u y   e s - v e   e t - e e   e u - e s   f a - i r   f i - f i   f o - f o   f r - b e   f r - c a   f r - c h   f r - f r   f r - l u   f r - m c   g l - e s   g u - i n   h e - i l   h i - i n   h r - b a   h r - h r   h u - h u   h y - a m   i d - i d   i s - i s   i t - c h   i t - i t   j a - j p   k a - g e   k k - k z   k n - i n   k o k - i n     k o - k r   k y - k g   l t - l t   l v - l v   m i - n z   m k - m k   m l - i n   m n - m n   m r - i n   m s - b n   m s - m y   m t - m t   n b - n o   n l - b e   n l - n l   n n - n o   n s - z a   p a - i n   p l - p l   p t - b r   p t - p t   q u z - b o     q u z - e c     q u z - p e     r o - r o   r u - r u   s a - i n   s e - f i   s e - n o   s e - s e   s k - s k   s l - s i   s m a - n o     s m a - s e     s m j - n o     s m j - s e     s m n - f i     s m s - f i     s q - a l   s r - b a - c y r l     s r - b a - l a t n     s r - s p - c y r l     s r - s p - l a t n     s v - f i   s v - s e   s w - k e   s y r - s y     t a - i n   t e - i n   t h - t h   t n - z a   t r - t r   t t - r u   u k - u a   u r - p k   u z - u z - c y r l     u z - u z - l a t n     v i - v n   x h - z a   z h - c h s     z h - c h t     z h - c n   z h - h k   z h - m o   z h - s g   z h - t w   z u - z a                     �      ���������������-DT�!�?-DT�!��RUUUUU�?        v�F�$I�?������ɿ��3Y�E�?#Y��q���n����?��;
9��� ��/I�?hK����d��?81�U����H!G�?��#�$�����0|f?�K�RVn���TUUUU�?        ~I�$I�?g����ɿHB�;E�?����q���{雮?�x��֚��                   �      �?       @       @      �?      �?      @>��1|�MC                     ���5�h!����?      �?            �?5�h!���>@�������             ��      �@      �                                                  �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������                                      �?1mm.�s�,�)���?   �'>�      �?�i����i<���?   �mb�      �?Z"�������.��?   ���u�      �?ϕk��|��c����}�?   ��,g�      �?y�sh:��;�8]+�?    �^<      �?ty�[g�ſ�h�9;��?    �%�<      �?���S�Ϳ�	%�L�?    jh<      �?2���y��?�;f���?    4݋�      �?Xw$��3�?Ak���?    �ł�      �?��暳s�?��)f��?   �0�9<      �?N��,J������8�?   ���v�      �?uZEeu��F�2�k��?    �Wt<      �?-��v1��?�-�VA��?   �`�<      �?�gY���\�ϗb�?    bu<      �?P/Ye���&%ѣ���?   @�}��      �?              �?                P/Ye��?&%ѣ���?   @�}��      ���gY�?�\�ϗb�?    bu<      п-��v1����-�VA��?   �`�<      пuZEeu�?F�2�k��?    �Wt<      �N��,J�?����8�?   ���v�      ࿇�暳s����)f��?   �0�9<      �Xw$��3��Ak���?    �ł�      �2���y�ʿ�;f���?    4݋�      ����S��?�	%�L�?    jh<      �ty�[g��?�h�9;��?    �%�<      �y�sh:�?;�8]+�?    �^<      �ϕk��|�?c����}�?   ��,g�      �Z"����?��.��?   ���u�      ��i��?�i<���?   �mb�      �1mm.�s?,�)���?   �'>�      �                              �1mm.�s?,�)����   �'><      ��i��?�i<��ȿ   �mb<      �Z"����?��.�ҿ   ���u<      �ϕk��|�?c����}ؿ   ��,g<      �y�sh:�?;�8]+޿    �^�      �ty�[g��?�h�9;��    �%��      ����S��?�	%�L�    jh�      �2���y�ʿ�;f���    4݋<      �Xw$��3��Ak���    �ł<      ࿇�暳s����)f��   �0�9�      �N��,J�?����8�   ���v<      �uZEeu�?F�2�k��    �Wt�      �-��v1����-�VA��   �`��      п�gY�?�\�ϗb�    bu�      пP/Ye��?&%ѣ���   @�}�<      ��              �                P/Ye���&%ѣ���   @�}�<      �?�gY���\�ϗb�    bu�      �?-��v1��?�-�VA��   �`��      �?uZEeu��F�2�k��    �Wt�      �?N��,J������8�   ���v<      �?��暳s�?��)f��   �0�9�      �?Xw$��3�?Ak���    �ł<      �?2���y��?�;f���    4݋<      �?���S�Ϳ�	%�L�    jh�      �?ty�[g�ſ�h�9;��    �%��      �?y�sh:��;�8]+޿    �^�      �?ϕk��|��c����}ؿ   ��,g<      �?Z"�������.�ҿ   ���u<      �?�i����i<��ȿ   �mb<      �?1mm.�s�,�)����   �'><      �?UUUUUUſ      ��?UUUUUU�?��*�l�l�V�4�V���>���>���m0_$@      8C  `a��=  `a��=  @T�!�?sp.�c;      `C      �<�������?       �      �?      ��������� �,�8�@�H�T�`�j��,�H�\�|�l�t�|������������������������������������������������������������� �������� �,�8�@�L�d�p����������$�H�d����������� ���<�D�P�`�|��������@�\���������j�__based(    __cdecl __pascal    __stdcall   __thiscall  __fastcall  __clrcall   __eabi  __ptr64 __restrict  __unaligned restrict(    new     delete =   >>  <<  !   ==  !=  []  operator    ->  *   ++  --  -   +   &   ->* /   %   <   <=  >   >=  ,   ()  ~   ^   |   &&  ||  *=  +=  -=  /=  %=  >>= <<= &=  |=  ^=  `vftable'   `vbtable'   `vcall' `typeof'    `local static guard'    `string'    `vbase destructor'  `vector deleting destructor'    `default constructor closure'   `scalar deleting destructor'    `vector constructor iterator'   `vector destructor iterator'    `vector vbase constructor iterator' `virtual displacement map'  `eh vector constructor iterator'    `eh vector destructor iterator' `eh vector vbase constructor iterator'  `copy constructor closure'  `udt returning' `EH `RTTI   `local vftable' `local vftable constructor closure'  new[]   delete[]   `omni callsig'  `placement delete closure'  `placement delete[] closure'    `managed vector constructor iterator'   `managed vector destructor iterator'    `eh vector copy constructor iterator'   `eh vector vbase copy constructor iterator' `dynamic initializer for '  `dynamic atexit destructor for '    `vector copy constructor iterator'  `vector vbase copy constructor iterator'    `managed vector copy constructor iterator'  `local static thread guard'  Type Descriptor'    Base Class Descriptor at (  Base Class Array'   Class Hierarchy Descriptor'     Complete Object Locator'   ������ �Sun Mon Tue Wed Thu Fri Sat Sunday  Monday  Tuesday Wednesday   Thursday    Friday  Saturday    Jan Feb Mar Apr May Jun Jul Aug Sep Oct Nov Dec January February    March   April   June    July    August  September   October November    December    AM  PM  MM/dd/yy    dddd, MMMM dd, yyyy HH:mm:ss    S u n   M o n   T u e   W e d   T h u   F r i   S a t   S u n d a y     M o n d a y     T u e s d a y   W e d n e s d a y   T h u r s d a y     F r i d a y     S a t u r d a y     J a n   F e b   M a r   A p r   M a y   J u n   J u l   A u g   S e p   O c t   N o v   D e c   J a n u a r y   F e b r u a r y     M a r c h   A p r i l   J u n e     J u l y     A u g u s t     S e p t e m b e r   O c t o b e r   N o v e m b e r     D e c e m b e r     A M     P M     M M / d d / y y     d d d d ,   M M M M   d d ,   y y y y   H H : m m : s s     (null)  ( n u l l )            EEE50 P    ( 8PX 700WP        `h````  xpxxxx              	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ 1#SNAN  1#IND   1#INF   1#QNAN                                                                                                                                                                                                                                                                                    ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������sinh    cosh    tanh    atan2   fabs    ldexp   _cabs   _hypot  fmod    frexp   _y0 _y1 _yn _logb   _nextafter  A      C O N O U T $   ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           � ��   RSDS��>��<L�VRVk   D:\Applications\MAXON\CINEMA 4D R14 Demo\plugins\AMa_1D_Snap\__build_win\obj\Win32_Release\AMa_1D_Snap_Win32_Release.pdb        �   �                  ���$�             ����    @   ��         ����    @   @�           P�$�               h�x��$�    0        ����    @   X�            T ��           ����x��$�    T        ����    @   ��             @�            l �            �(�    l         ����    @   �            � X�           h�p�    �         ����    @   X�    �� ��                      ����    ����    ����    ˎ    ����    ����    ����c�}�    ����    ����    ����    ʘ    ����    ����    ����    ��    ����    ����    ����    ������    ������    ����    ����    �����    .�����    ����    ����    ��    ����    |���    ����    k�    ����    ����    ����    W�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    2�    ����    ����    ����    ��    ����    ����    ����y���    ����    ����    ������    ����    ����    ����    Y    ����    ����    ����    	<        �;����    ����    ����    �<    ����    ����    ����    h=    ����    ����    ����    �F    ����    ����    ����9NUN    ����    ����    ����    �Q    ����    ����    ����    �R    ����    ����    ����    GS    ����    ����    ����    W�         ��  `                     �  � 0� B� X� h� t� �� �� �� �� �� �� �� � � 2� D� Z� l� z� �� �� �� �� �� � ,� F� `� v� �� �� �� �� �� ��  � 
� � &� :� F� \� n� ~� �� �� �� �� �� �� �� �� � � .� @� T� f� z� �� �� ��     <EncodePointer DecodePointer �GetCommandLineA (GetCurrentThreadId  jGetLastError  QHeapFree  MHeapAlloc �GetStdHandle  �WriteFile }GetModuleFileNameW  �IsProcessorFeaturePresent SetLastError  qInterlockedIncrement  mInterlockedDecrement  mExitProcess �GetModuleHandleExW  �GetProcAddress  �MultiByteToWideChar �GetProcessHeap  WGetFileType fInitializeCriticalSectionAndSpinCount DeleteCriticalSection �GetStartupInfoW |GetModuleFileNameA  <QueryPerformanceCounter $GetCurrentProcessId �GetSystemTimeAsFileTime @GetEnvironmentStringsW  �FreeEnvironmentStringsW �WideCharToMultiByte �UnhandledExceptionFilter  PSetUnhandledExceptionFilter #GetCurrentProcess oTerminateProcess  �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree �GetModuleHandleW  _Sleep �IsDebuggerPresent VHeapSize  OutputDebugStringW  �LoadLibraryExW  �LoadLibraryW  �LCMapStringW  @EnterCriticalSection  �LeaveCriticalSection  �RtlUnwind �IsValidCodePage �GetACP  �GetOEMCP  �GetCPInfo THeapReAlloc �GetStringTypeW  �GetConsoleCP  GetConsoleMode  	SetFilePointerEx  HRaiseException  �FlushFileBuffers  /SetStdHandle  �WriteConsoleW � CloseHandle � CreateFileW KERNEL32.dll                  `�
R    �          �� ��  � P� �   AMa_1D_Snap.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      dz    .?AVToolData@@  dz    .?AVBaseData@@  dz    .?AVDescriptionToolData@@   dz    .?AVD1Snap@@    dz    .?AVNeighbor@@              dz    .?AVtype_info@@ u�  s�  N�@���D                       atan            cos             sin             ������������������������    �����
                                                          ����                                             	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                sqrt            �&                                                                                                                                                                                                                                                                                                @�  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                                                                                                                                                                                                                                                                                                   abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                                     abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                            C       ���������������������������������� �$�(�,�0�4�8�@�L�T��\�d�l�t�����������������       ���������������,�<�P�d�t���������������������������������$�0�<�L�`�p�������������<��
                                   `	            `	            `	            `	            `	                          8        ����h	                           ���� !     !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �� �         �            8.   4 ! ! ! ! ! ! ! ! !�!!!!!!!.   �   ���5      @   �  �   ����             ��           D�   H�   8�   <�   �    �!   (�   L�   T�   d�   0�   ��   ��   ��    ��   l�   t�   8�   |�   @�   H�   P�   X�   `�"   h�#   l�$   p�%   t�&   |�       �D        � 0                  �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
          �      ���������              �����                                                                                                                                                                                                                                                                                                                               �   
0�0�2�2�233k3�35C5_5�5�5�5606d6�6p7x7J8R8$9,9�9:t:�:�:;�;�;�;�;<1<9<A<I<a<�<�<�<�<�<�=�=>>5>L>b>y>�>�>�>?*?:?l?~?�?�?    p   0[0`0�0�0�0�1<2�2�3�3464I4�4�4�4�4�4�45Q5y5�546X637a7{7�7�7�7	8*8Y8�8�89"9u:�:�<�<"=�=>Q>i>�>�>�?   0  �   00<0b0|0�0�0�01x1|1�1�1�1�1�1�1=2p2�2�2�2�2�233�3�5�5f6�6W7�7�7 8D8]8y8�8�8�8�8�89D9^9u9�9�9|:�:�:;�;�;<5<�<�<F='>;>P>a>w>�>�>�>�>�>??A?X?s?�?�?�?�?�? @  0   0070N0y0�0�0�0�0�021�1}2�25�6�8=�>   P  (   �3�5�:;U;�;�;R<y<�<�<�<�<=D=Q> `  �   �0�0�0�0141a1�1�1�1�1%232A2V2h2z2�2�2�2�2�2�2�23*3;3L3�3�34N4�4�4�4�4�4	55/5u5�5�5�5�5�56%6�6�6�6�67%7�7�7	8%8�8�8�8�89.9T9�9�9�9+:G:�:�:�:F;e;�;<y<�<�<�<�<==$=a=t=�=�=�=�=>!>4>T>|>�>�>�>??D?d?�?�?�?�?�? p  �   040Q0t0�1�1�1�1�1�1�1�1�1�1�1 22222#2�2�2�2h3�34D4Z4�4�4�455A5T5�5�5�56!6A6g6�6�6�6717Q7q7�7�7�78$8D8d8�8�8�8�89!949T9t9�9�9�9�9�:�:";�;�;V<w<�<=7=�=+>B>�>P?j?�?   �  �   ]0w0�0�0�0L1�1�12 2W2�2�2$3�3�3�34G4�4-5G5d5�5�56�6�617�7�7�7 878�8 9:9�90:J:�:;!;G;t;�;�;�;<8<s<�<�<�<==2=O=]=�=�=�=>!>D>a>t>�>�>�>?G?w?�?�?�?�?   �  �   040T0t0�0�0�0�0�0�0�0!111D1d1�1�1�1�1242d2�2�2�2+3c3�3�334t4�4�4�4q5�5�5�5�5'6Q6d6�6�6�67'7T7w7�7�7�7$8G8�8�8�8�8�8�89$9A9Q9d9�9�9�9�9:4:H:Z:b:s:�:�:�:�:�:�:;4;N;b;r;�;�;�;�;�;<4<T<t<�<�<�<�<=!=1=D=d=�=�=�=�=>0>T>t>�>�>�>�>?$?D?�?�?�? �  �   040T0t0�0�0�0�01$1D1d1�1�1�1�1�122%2D2d2�2�23D3d3�3�3�3�34$4D4�4�4�4�4�4,515M5b5�5�56Q6t6�6�6�6!747d7�7�7�78*8H8m8�8�8�8�89<9P9`9�9�9�9�9:4:L:l:�:�:�:�:;-;M;t;�;�;�;�;�;<5<M<m<�<�<�<�<�<===U=u=�=�=�=�=>5>U>|>�>�>�>�>?>?d?�?�?�?�? �  �   0!040T0t0�0�0�0�0�0$1D1d1�1�1�1�12$2D2d2�2�2�2�2�23$3L3g3�3�3�3'4W4�4�4�4Y5'6T6q6�6�6�6�6777d7�7�7�7�7'8W8�8�8�89'9\9�9�9�9:4:Q:t:�:�:�:�:;D;q;�;�;<D<t<�<�<�<0=O=g=�=�=�=>!>D>T>�>�>�>�>$?;?e?�?�?�?   �  �   00:0\0o0�0�0�0111Q1q1�1�1�1!2D2d2�2�2�23G3q3�3�3�34$4D4t4�4�4
555I5g5�5�5�5�5616T6�6�6�677u7�78w8�8�8�8949V9{9�9�9�9A:d:�:�:�:;$;A;d;�;�;�;�;<D<d<�<�<�<�<=7=d=�=�=�=�=>$>A>q>�>�>?a?�?�?�?   �  �   0?0|0�0�01H1w1�1�1�1�1262M243?3�3�3�3�3�3B4B6�8�8=9E9~9�9�9�9:�;�;�;�;�;<$<L<�<�<�<=%=*=D=l=�=�=>4>W>�>�>K?�?�?�?�?   �  �   70q0�0�0�0�1�1�4�4�4545Q5t5�5�5�56$6D6a6�6�6�67o7�788p8�8�839k9�9�9 :E:J:u:�:�:�:�:�:�:�:�:;(;B;m;�;�;�;�;�;�;<<*<;<M<U<t<�<�<�<�<�<
==1=E=e==�=�=�=�=�=�=>>+>=>E>d>x>�>�>�>�>�>?!?5?U?o?�?�?�?�?�?�?   �    00+0U0d0p0�0�0�0�0�0�0�01!1M1g1x1�1�1�1�1�1�12"2*2I2]2}2�2�2�2�2�2�23/3@3S3x3�344>4�4�4�4�4�45<5P5p5�5�5�5�5�5U6f6w66�6�67757I7[7l7�7�7�7�718B8K8T8f8q8�8�8�89A9g9�9�9�9:4:d:�:�:b;k;r;y;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<G<t<�<>$>_>�>�>�>i?�?   �   d0�01�1:2�2�2�2�2!3�34�4b5�5�5�56u6�6�6�6!7U7}7�7�7858u8�8�89%9e9�9�91:b:�:�:�:;Q;y;�;�;�;�;<,<Q<y<�<�<=W=�=�=�=->m>�>�>2?b?�?�?  �   0R0�0�01U1�1�12E2u2�2�253�3�3�3%4V4�4�4%5e5�5�5%6u6�67D7x7�7�7�7�78'818D8g8�8�8�8�8�899#9D9U9c9�9�9�9�9�9:,:@:P:t:�:�:�:�:�:�:;,;@;N;];o;�;�;�;�;�;�;!<1<D<d<�<�<�<�<=!=4=d=v=�=�=�=�=>$><>P>`>�>�>�>�>�>?7?Q?a?q?�?�?�?�?       0$0D0d0�0�0�0�01.1U1�1�1�1�12#2m2�2�2�23343d3�3�3�3�3�344R4m4�4�4�45$5D5d5�5�5�5�5646T6p6�6�6�6�677!7<7p7�7�7�78D8h8�8�8�89.9P9r9�9�9�9:<:`:�:�:�:!;4;d;�;�;�;�;<<!<1<A<Q<d<�<�<�<�<�<�<=$=Q=a=t=�=�=�=�=�=�=>">2>Q>d>�>�>�>�>?4?T?t?�?�?�?�?   0   0D0d0�0�0�0�0141T1t1�1�1�1�1242a2�2�2�2�23$3D3d3�3�3�3�34$4D4d4�4�4�4�45$5D5d5�5�5�5�5616D6d6�6�6�6�6�677!717D7t7�7�7�7�7�7848T8t8�8�8�899=9O9t9�9�9�9�9:4:K:_:m:|:�:�:�:�:�:�:;X;};�;�;�;�;�;�;<<D<a<u<�<�<�<�<�<=$=D=X=h=�=�=�=�=>D>d>�>�>�>?D?d?�?�?�?�?�? @ �   040Q0a0q0�0�0�0�0111W1�1�1�1�1�1272g2�2�2�23T3g3{3�3�34!4A4a4�4�4�4�45F5Y5�5�5�5�516F6P6�677l7�7�7�7818D8�9�9�9:y:~:;G<t<�<�<�<�<�>�>?-?�?   P �   0~1�1�1�2�2�2�2343T3q3�3�3�3�34$4A4q4�4�4�45<5t5�5�5�5�56!646T6t6�6�6�6�6�67!717D7d7�7�7�7�78.8Q8d8�8�8�8�899D9u9�9�9�9�9�9:Q:t:�:�:�:;!;D;T;�;�;�;�;<$<Q<q<�<�<�<�<=4=T=�=�=�=�=>1>T>t>�>�>D?�?�?�?   ` h   040T0t0�0�0�01$1A1d1�1�1�172a2�2O3T3u3z3�3�344�4575<566=6B6�6767;7�7�7�9:N?�?�?�?�?�?   p T   <2�2�2�518]8�8�89U9�9�9:B:u:�:�:%;e;�;�;"<R<�<�<�<=U=�=�=>U>�>�>?e?�?   �   0U0�0�0%1�1�2�2�23>3a3�3d4q4w4�4�4�455-5D5H5L5P5T5X5l5t5�5�546d6�6�6�67767B7N7Z77�7�7�7�7�7�7�7�78(808Q8e8�8�8�8�8�8�8�89969J9c9l9::(:4:Q:W:l:�:�:�:R;�;�;�;�;<<,<Q<�<�<=='=K=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�='>,>6>j>>�>�>�>�>?.?�?�?�?   �    0D0�0�0�0�0111@1�1�12C2k2y2%4C4\4c4k4p4t4x4�4�4�4�4�4�4�4�4 555R5X5\5`5d5�5�5�5�5�5 66%6O6�6�6�6�6�6�6�6�6�6�6�6�6�6 7u8z88�8�8�8�8Z9_9h9t9y9�9�9�9�;�;�;�;�;�;�;�;!<G<e<l<p<t<x<|<�<�<�<�<�<�<�<�<J=U=p=w=|=�=�=�=�=>>>>>>> >$>n>t>x>|>�> � �   141G1W1�1�1�1�1�1�1�1�1
22'2.272P2Z2�2�2�23R3h3p3v33�3(4a4j4y4�4�4�4�4�4�4�4'5A5H5Q5Z5c5l5x5�5�5�5�5�5666666 6$6(6,6064686<6B6�6�6�67'7=7O7b7�7	88)848a8l8~8�8�899G9Y9d9�9�9�9O:p:u:�:�:;; � �   "0y0�0p2/3�56	6�7888B8z8�8�8�899H9c9{9�9�9�9�9�9N:Y:z:�:�:�:�:�:�:�:;;;";@;M;V;q;};�;�;�;�;�;�;�;�;�;�;�;�;�;<
<<R<Z<m<x<}<�<�<�<�<�<�<�<}=�=�=�=�=�=�=�=	>>>$>G>L>X>]>|>�>�>�>�>�>??O?[?�?�?�? � �  0&0I0O0V0�0�0�0&1?1w1�1�1�1�1�1�1�1�1a2g2�34=4G4�4�4�4�4�4�4�4
55"5/5^5f5u5�5�5�5�5�5666!606:6@6O6Y6_6q6~6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�67777 7%7+73787>7F7K7Q7Y7^7d7l7q7w77�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78	8888"8*8/858=8B8H8P8U8[8c8h8n8v8{8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8999>9G9U9q9�9�9�9�9�9::!:&:A:^:�:L;T;k;�;�;?<s<�<�<�<�<�<�=�=�=�=>>!>3>=>_>j>�>�?�?�? � ,  0000%0+02090@0G0N0U0\0d0l0t0�0�0�0�0�0�0�0�0�0�011`1r1�1�1�1�1�2333�5�5�5�5�56$6*666D6J6Y6`6p6v6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6777!7d7|7�7�7�7�7�7�7�7�73888w8|8�8�8�8�8�899)939�9:9:b:p:v:�:1;j;r;�;�;�;�;�;�;�;<(<4<@<L<X<d<p<�<�<�<�<�<== =8=D=P=\=�=�=�=�=�=�=�=�=�=Y>�>h?�?   � �   ;0<1L1]1e1u1�1)252E2Q2n2t2�2�2�2�2~3�3�3�344$494^4�4�4*5@5P5�5�5�5�5
6636<6H6S6x6�6�6�6�6�677*707U7a7l8�8�889�9%:�:�:;,;e;�;�;�;<"<)<0<K<W<a<n<x<�<�<=0=�>�>�>�>�>?? ?A?�?�?�?�?   � �   00"090S0n0w0}0�0�0�0�0�0�0-1c1v12C2j2�263A3�4�4�6J7�8�:�:;+;?;E;�;<<!<-<4<N<]<j<v<�<�<�<�<�<�<�<�<�<=<=I=R=v=�=N>T>`>�>�>�>??     P   +020�041;1a1h1�1�12r5_6�7�7�78$8*8�9�;�;�;�;�;<<<�<X=>�>a?m?�?�?    h   0;0M0_0q0�0�0�0�0�0�0�01121D1V1h1z15u5�5�6<7y7�7899#979C9�9':I;Q;�<�=�=%>+>9>H>�>�> ?�?     L   �0�0i2�23�3�3�3�3D4[4�45n8�8�;�;�;�;�;�;�;�;�;�;�;<<�<�<�<=w=�= 0 <   �7K:\:7;];h;�;�;<<<C<j<w<|<�<�<�<=!=�=>�>�>�>�>I? @ `   050>0�0�0q1}1�1e2n2`3i3U4�4�4�4#575~5�5 66<6�6 7737v7�7_8{8�9�9�9�9�9%=>>(>Z>�>�>�> P h   1,1I1i1~1�1S2�2�23.3:3a3q3�3�3�3�34T4`4�4.5v5�5�5�67,7H7�7 8
8&8y8�8�8�8�8�8�8�8�8�8�8�899 ` T   1111 1$1014181�1�1�1�1�1�1 22222222 2$2(2,2024282<2@2D2�3�3�4�4�4 p    `:d:h:   � 8   �23333$3,343<3D3L3T3\3d3l3t3|3�3�3�3�3�3�3   � �  �0 1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12222$2,242<2D2L2T2\2d2l2t2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23333$3,343<3D3L3T3\3d3l3t3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�34444$4,444<4D4L4T4\4d4l4t4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�45555$5,545<5D5L5T5\5d5l5t5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�56666$6,646<6D6L6T6\6d6l6t6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�67777$7,747<7D7L7T7\7d7l7t7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78888$8,848<8D8L8T8\8d8l8t8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 9999 9(90989@9H9P9X9`9h9p9x9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::: :(:0:8:@:H:P:X:`:h:p:x:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;; ;(;0;8;@;H;P;X;`;h;p;x;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<< <(<0<8<@<H<P<X<`<h<p<x<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ==== =(=0=8=@=H=P=X=`=h=p=x=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>> >(>0>8>@>H>P>X>`>h>p>x>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???? ?(?0?8?@?H?P?X?`?h?p?x?�?�?�?�?�?�?�?�? � �   `5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�<�<�<�< � �   <:@:�:�: ;; ;$;<;L;P;d;h;l;p;x;�;�;�;�;�;�;�;�;�;�;�;�;<<< <(<@<P<T<d<h<p<�<�<�<�<=(=H=T=p=|=�=�=�=�=>8>X>t>x>�>�>�>�>�> ? ?@?\?`?�?�?�?�?   \   0000T0l0�0 11111111 1$1@4h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;$;4;T;`;d;h;l;�;�;>>0>8><>@>D>H>L>P>T>X>\>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>????$?,?4?<?D?L?T?\?d?l?t?|?�?�?�?�?�?�?�?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                